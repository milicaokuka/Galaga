
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 14			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

-- GENERATED BY BC_MEM_PACKER
-- DATE: Mon Jun 06 17:39:44 2016

	signal mem : ram_t := (

--	***** COLOR PALLETE *****


		
		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00DE6800", -- R: 0 G: 104 B: 222
		2 =>	x"00DEDEDE", -- R: 222 G: 222 B: 222
		3 =>	x"000000FF", -- R: 255 G: 0 B: 0
		4 =>	x"00DEB8B8", -- R: 184 G: 184 B: 222
		5 =>	x"00BCBCBC", -- R: 188 G: 188 B: 188
		6 =>	x"000028D8", -- R: 216 G: 40 B: 0
		7 =>	x"00EC3820", -- R: 32 G: 56 B: 236
		8 =>	x"00FCFCFC", -- R: 252 G: 252 B: 252
		9 =>	x"00DE00FF", -- R: 255 G: 0 B: 222
		10 =>	x"00DE0097", -- R: 151 G: 0 B: 222
		11 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		12 =>	x"00979700", -- R: 0 G: 151 B: 151
		13 =>	x"000047DE", -- R: 222 G: 71 B: 0
		14 =>	x"00000000", -- R: 0 G: 0 B: 0
		15 =>	x"00000000", -- R: 0 G: 0 B: 0
		16 =>	x"00000000", -- R: 0 G: 0 B: 0
		17 =>	x"00000000", -- R: 0 G: 0 B: 0
		18 =>	x"00000000", -- R: 0 G: 0 B: 0
		19 =>	x"00000000", -- R: 0 G: 0 B: 0
		20 =>	x"00000000", -- R: 0 G: 0 B: 0
		21 =>	x"00000000", -- R: 0 G: 0 B: 0
		22 =>	x"00000000", -- R: 0 G: 0 B: 0
		23 =>	x"00000000", -- R: 0 G: 0 B: 0
		24 =>	x"00000000", -- R: 0 G: 0 B: 0
		25 =>	x"00000000", -- R: 0 G: 0 B: 0
		26 =>	x"00000000", -- R: 0 G: 0 B: 0
		27 =>	x"00000000", -- R: 0 G: 0 B: 0
		28 =>	x"00000000", -- R: 0 G: 0 B: 0
		29 =>	x"00000000", -- R: 0 G: 0 B: 0
		30 =>	x"00000000", -- R: 0 G: 0 B: 0
		31 =>	x"00000000", -- R: 0 G: 0 B: 0
		32 =>	x"00000000", -- R: 0 G: 0 B: 0
		33 =>	x"00000000", -- R: 0 G: 0 B: 0
		34 =>	x"00000000", -- R: 0 G: 0 B: 0
		35 =>	x"00000000", -- R: 0 G: 0 B: 0
		36 =>	x"00000000", -- R: 0 G: 0 B: 0
		37 =>	x"00000000", -- R: 0 G: 0 B: 0
		38 =>	x"00000000", -- R: 0 G: 0 B: 0
		39 =>	x"00000000", -- R: 0 G: 0 B: 0
		40 =>	x"00000000", -- R: 0 G: 0 B: 0
		41 =>	x"00000000", -- R: 0 G: 0 B: 0
		42 =>	x"00000000", -- R: 0 G: 0 B: 0
		43 =>	x"00000000", -- R: 0 G: 0 B: 0
		44 =>	x"00000000", -- R: 0 G: 0 B: 0
		45 =>	x"00000000", -- R: 0 G: 0 B: 0
		46 =>	x"00000000", -- R: 0 G: 0 B: 0
		47 =>	x"00000000", -- R: 0 G: 0 B: 0
		48 =>	x"00000000", -- R: 0 G: 0 B: 0
		49 =>	x"00000000", -- R: 0 G: 0 B: 0
		50 =>	x"00000000", -- R: 0 G: 0 B: 0
		51 =>	x"00000000", -- R: 0 G: 0 B: 0
		52 =>	x"00000000", -- R: 0 G: 0 B: 0
		53 =>	x"00000000", -- R: 0 G: 0 B: 0
		54 =>	x"00000000", -- R: 0 G: 0 B: 0
		55 =>	x"00000000", -- R: 0 G: 0 B: 0
		56 =>	x"00000000", -- R: 0 G: 0 B: 0
		57 =>	x"00000000", -- R: 0 G: 0 B: 0
		58 =>	x"00000000", -- R: 0 G: 0 B: 0
		59 =>	x"00000000", -- R: 0 G: 0 B: 0
		60 =>	x"00000000", -- R: 0 G: 0 B: 0
		61 =>	x"00000000", -- R: 0 G: 0 B: 0
		62 =>	x"00000000", -- R: 0 G: 0 B: 0
		63 =>	x"00000000", -- R: 0 G: 0 B: 0
		64 =>	x"00000000", -- R: 0 G: 0 B: 0
		65 =>	x"00000000", -- R: 0 G: 0 B: 0
		66 =>	x"00000000", -- R: 0 G: 0 B: 0
		67 =>	x"00000000", -- R: 0 G: 0 B: 0
		68 =>	x"00000000", -- R: 0 G: 0 B: 0
		69 =>	x"00000000", -- R: 0 G: 0 B: 0
		70 =>	x"00000000", -- R: 0 G: 0 B: 0
		71 =>	x"00000000", -- R: 0 G: 0 B: 0
		72 =>	x"00000000", -- R: 0 G: 0 B: 0
		73 =>	x"00000000", -- R: 0 G: 0 B: 0
		74 =>	x"00000000", -- R: 0 G: 0 B: 0
		75 =>	x"00000000", -- R: 0 G: 0 B: 0
		76 =>	x"00000000", -- R: 0 G: 0 B: 0
		77 =>	x"00000000", -- R: 0 G: 0 B: 0
		78 =>	x"00000000", -- R: 0 G: 0 B: 0
		79 =>	x"00000000", -- R: 0 G: 0 B: 0
		80 =>	x"00000000", -- R: 0 G: 0 B: 0
		81 =>	x"00000000", -- R: 0 G: 0 B: 0
		82 =>	x"00000000", -- R: 0 G: 0 B: 0
		83 =>	x"00000000", -- R: 0 G: 0 B: 0
		84 =>	x"00000000", -- R: 0 G: 0 B: 0
		85 =>	x"00000000", -- R: 0 G: 0 B: 0
		86 =>	x"00000000", -- R: 0 G: 0 B: 0
		87 =>	x"00000000", -- R: 0 G: 0 B: 0
		88 =>	x"00000000", -- R: 0 G: 0 B: 0
		89 =>	x"00000000", -- R: 0 G: 0 B: 0
		90 =>	x"00000000", -- R: 0 G: 0 B: 0
		91 =>	x"00000000", -- R: 0 G: 0 B: 0
		92 =>	x"00000000", -- R: 0 G: 0 B: 0
		93 =>	x"00000000", -- R: 0 G: 0 B: 0
		94 =>	x"00000000", -- R: 0 G: 0 B: 0
		95 =>	x"00000000", -- R: 0 G: 0 B: 0
		96 =>	x"00000000", -- R: 0 G: 0 B: 0
		97 =>	x"00000000", -- R: 0 G: 0 B: 0
		98 =>	x"00000000", -- R: 0 G: 0 B: 0
		99 =>	x"00000000", -- R: 0 G: 0 B: 0
		100 =>	x"00000000", -- R: 0 G: 0 B: 0
		101 =>	x"00000000", -- R: 0 G: 0 B: 0
		102 =>	x"00000000", -- R: 0 G: 0 B: 0
		103 =>	x"00000000", -- R: 0 G: 0 B: 0
		104 =>	x"00000000", -- R: 0 G: 0 B: 0
		105 =>	x"00000000", -- R: 0 G: 0 B: 0
		106 =>	x"00000000", -- R: 0 G: 0 B: 0
		107 =>	x"00000000", -- R: 0 G: 0 B: 0
		108 =>	x"00000000", -- R: 0 G: 0 B: 0
		109 =>	x"00000000", -- R: 0 G: 0 B: 0
		110 =>	x"00000000", -- R: 0 G: 0 B: 0
		111 =>	x"00000000", -- R: 0 G: 0 B: 0
		112 =>	x"00000000", -- R: 0 G: 0 B: 0
		113 =>	x"00000000", -- R: 0 G: 0 B: 0
		114 =>	x"00000000", -- R: 0 G: 0 B: 0
		115 =>	x"00000000", -- R: 0 G: 0 B: 0
		116 =>	x"00000000", -- R: 0 G: 0 B: 0
		117 =>	x"00000000", -- R: 0 G: 0 B: 0
		118 =>	x"00000000", -- R: 0 G: 0 B: 0
		119 =>	x"00000000", -- R: 0 G: 0 B: 0
		120 =>	x"00000000", -- R: 0 G: 0 B: 0
		121 =>	x"00000000", -- R: 0 G: 0 B: 0
		122 =>	x"00000000", -- R: 0 G: 0 B: 0
		123 =>	x"00000000", -- R: 0 G: 0 B: 0
		124 =>	x"00000000", -- R: 0 G: 0 B: 0
		125 =>	x"00000000", -- R: 0 G: 0 B: 0
		126 =>	x"00000000", -- R: 0 G: 0 B: 0
		127 =>	x"00000000", -- R: 0 G: 0 B: 0
		128 =>	x"00000000", -- R: 0 G: 0 B: 0
		129 =>	x"00000000", -- R: 0 G: 0 B: 0
		130 =>	x"00000000", -- R: 0 G: 0 B: 0
		131 =>	x"00000000", -- R: 0 G: 0 B: 0
		132 =>	x"00000000", -- R: 0 G: 0 B: 0
		133 =>	x"00000000", -- R: 0 G: 0 B: 0
		134 =>	x"00000000", -- R: 0 G: 0 B: 0
		135 =>	x"00000000", -- R: 0 G: 0 B: 0
		136 =>	x"00000000", -- R: 0 G: 0 B: 0
		137 =>	x"00000000", -- R: 0 G: 0 B: 0
		138 =>	x"00000000", -- R: 0 G: 0 B: 0
		139 =>	x"00000000", -- R: 0 G: 0 B: 0
		140 =>	x"00000000", -- R: 0 G: 0 B: 0
		141 =>	x"00000000", -- R: 0 G: 0 B: 0
		142 =>	x"00000000", -- R: 0 G: 0 B: 0
		143 =>	x"00000000", -- R: 0 G: 0 B: 0
		144 =>	x"00000000", -- R: 0 G: 0 B: 0
		145 =>	x"00000000", -- R: 0 G: 0 B: 0
		146 =>	x"00000000", -- R: 0 G: 0 B: 0
		147 =>	x"00000000", -- R: 0 G: 0 B: 0
		148 =>	x"00000000", -- R: 0 G: 0 B: 0
		149 =>	x"00000000", -- R: 0 G: 0 B: 0
		150 =>	x"00000000", -- R: 0 G: 0 B: 0
		151 =>	x"00000000", -- R: 0 G: 0 B: 0
		152 =>	x"00000000", -- R: 0 G: 0 B: 0
		153 =>	x"00000000", -- R: 0 G: 0 B: 0
		154 =>	x"00000000", -- R: 0 G: 0 B: 0
		155 =>	x"00000000", -- R: 0 G: 0 B: 0
		156 =>	x"00000000", -- R: 0 G: 0 B: 0
		157 =>	x"00000000", -- R: 0 G: 0 B: 0
		158 =>	x"00000000", -- R: 0 G: 0 B: 0
		159 =>	x"00000000", -- R: 0 G: 0 B: 0
		160 =>	x"00000000", -- R: 0 G: 0 B: 0
		161 =>	x"00000000", -- R: 0 G: 0 B: 0
		162 =>	x"00000000", -- R: 0 G: 0 B: 0
		163 =>	x"00000000", -- R: 0 G: 0 B: 0
		164 =>	x"00000000", -- R: 0 G: 0 B: 0
		165 =>	x"00000000", -- R: 0 G: 0 B: 0
		166 =>	x"00000000", -- R: 0 G: 0 B: 0
		167 =>	x"00000000", -- R: 0 G: 0 B: 0
		168 =>	x"00000000", -- R: 0 G: 0 B: 0
		169 =>	x"00000000", -- R: 0 G: 0 B: 0
		170 =>	x"00000000", -- R: 0 G: 0 B: 0
		171 =>	x"00000000", -- R: 0 G: 0 B: 0
		172 =>	x"00000000", -- R: 0 G: 0 B: 0
		173 =>	x"00000000", -- R: 0 G: 0 B: 0
		174 =>	x"00000000", -- R: 0 G: 0 B: 0
		175 =>	x"00000000", -- R: 0 G: 0 B: 0
		176 =>	x"00000000", -- R: 0 G: 0 B: 0
		177 =>	x"00000000", -- R: 0 G: 0 B: 0
		178 =>	x"00000000", -- R: 0 G: 0 B: 0
		179 =>	x"00000000", -- R: 0 G: 0 B: 0
		180 =>	x"00000000", -- R: 0 G: 0 B: 0
		181 =>	x"00000000", -- R: 0 G: 0 B: 0
		182 =>	x"00000000", -- R: 0 G: 0 B: 0
		183 =>	x"00000000", -- R: 0 G: 0 B: 0
		184 =>	x"00000000", -- R: 0 G: 0 B: 0
		185 =>	x"00000000", -- R: 0 G: 0 B: 0
		186 =>	x"00000000", -- R: 0 G: 0 B: 0
		187 =>	x"00000000", -- R: 0 G: 0 B: 0
		188 =>	x"00000000", -- R: 0 G: 0 B: 0
		189 =>	x"00000000", -- R: 0 G: 0 B: 0
		190 =>	x"00000000", -- R: 0 G: 0 B: 0
		191 =>	x"00000000", -- R: 0 G: 0 B: 0
		192 =>	x"00000000", -- R: 0 G: 0 B: 0
		193 =>	x"00000000", -- R: 0 G: 0 B: 0
		194 =>	x"00000000", -- R: 0 G: 0 B: 0
		195 =>	x"00000000", -- R: 0 G: 0 B: 0
		196 =>	x"00000000", -- R: 0 G: 0 B: 0
		197 =>	x"00000000", -- R: 0 G: 0 B: 0
		198 =>	x"00000000", -- R: 0 G: 0 B: 0
		199 =>	x"00000000", -- R: 0 G: 0 B: 0
		200 =>	x"00000000", -- R: 0 G: 0 B: 0
		201 =>	x"00000000", -- R: 0 G: 0 B: 0
		202 =>	x"00000000", -- R: 0 G: 0 B: 0
		203 =>	x"00000000", -- R: 0 G: 0 B: 0
		204 =>	x"00000000", -- R: 0 G: 0 B: 0
		205 =>	x"00000000", -- R: 0 G: 0 B: 0
		206 =>	x"00000000", -- R: 0 G: 0 B: 0
		207 =>	x"00000000", -- R: 0 G: 0 B: 0
		208 =>	x"00000000", -- R: 0 G: 0 B: 0
		209 =>	x"00000000", -- R: 0 G: 0 B: 0
		210 =>	x"00000000", -- R: 0 G: 0 B: 0
		211 =>	x"00000000", -- R: 0 G: 0 B: 0
		212 =>	x"00000000", -- R: 0 G: 0 B: 0
		213 =>	x"00000000", -- R: 0 G: 0 B: 0
		214 =>	x"00000000", -- R: 0 G: 0 B: 0
		215 =>	x"00000000", -- R: 0 G: 0 B: 0
		216 =>	x"00000000", -- R: 0 G: 0 B: 0
		217 =>	x"00000000", -- R: 0 G: 0 B: 0
		218 =>	x"00000000", -- R: 0 G: 0 B: 0
		219 =>	x"00000000", -- R: 0 G: 0 B: 0
		220 =>	x"00000000", -- R: 0 G: 0 B: 0
		221 =>	x"00000000", -- R: 0 G: 0 B: 0
		222 =>	x"00000000", -- R: 0 G: 0 B: 0
		223 =>	x"00000000", -- R: 0 G: 0 B: 0
		224 =>	x"00000000", -- R: 0 G: 0 B: 0
		225 =>	x"00000000", -- R: 0 G: 0 B: 0
		226 =>	x"00000000", -- R: 0 G: 0 B: 0
		227 =>	x"00000000", -- R: 0 G: 0 B: 0
		228 =>	x"00000000", -- R: 0 G: 0 B: 0
		229 =>	x"00000000", -- R: 0 G: 0 B: 0
		230 =>	x"00000000", -- R: 0 G: 0 B: 0
		231 =>	x"00000000", -- R: 0 G: 0 B: 0
		232 =>	x"00000000", -- R: 0 G: 0 B: 0
		233 =>	x"00000000", -- R: 0 G: 0 B: 0
		234 =>	x"00000000", -- R: 0 G: 0 B: 0
		235 =>	x"00000000", -- R: 0 G: 0 B: 0
		236 =>	x"00000000", -- R: 0 G: 0 B: 0
		237 =>	x"00000000", -- R: 0 G: 0 B: 0
		238 =>	x"00000000", -- R: 0 G: 0 B: 0
		239 =>	x"00000000", -- R: 0 G: 0 B: 0
		240 =>	x"00000000", -- R: 0 G: 0 B: 0
		241 =>	x"00000000", -- R: 0 G: 0 B: 0
		242 =>	x"00000000", -- R: 0 G: 0 B: 0
		243 =>	x"00000000", -- R: 0 G: 0 B: 0
		244 =>	x"00000000", -- R: 0 G: 0 B: 0
		245 =>	x"00000000", -- R: 0 G: 0 B: 0
		246 =>	x"00000000", -- R: 0 G: 0 B: 0
		247 =>	x"00000000", -- R: 0 G: 0 B: 0
		248 =>	x"00000000", -- R: 0 G: 0 B: 0
		249 =>	x"00000000", -- R: 0 G: 0 B: 0
		250 =>	x"00000000", -- R: 0 G: 0 B: 0
		251 =>	x"00000000", -- R: 0 G: 0 B: 0
		252 =>	x"00000000", -- R: 0 G: 0 B: 0
		253 =>	x"00000000", -- R: 0 G: 0 B: 0
		254 =>	x"00000000", -- R: 0 G: 0 B: 0
		

		
		
--			***** 8x8 IMAGES *****




--		***** 16x16 IMAGES *****


		-- GENERATED BY BC_MEM_PACKER
-- DATE: Fri May 19 14:46:42 2017



--			***** 8x8 IMAGES *****




--			***** 16x16 IMAGES *****


		255 =>	x"00000000", -- IMG_16x16_avion2_10
		256 =>	x"00010000",
		257 =>	x"00000000",
		258 =>	x"00000000",
		259 =>	x"00000101",
		260 =>	x"01010100",
		261 =>	x"00020100",
		262 =>	x"00000000",
		263 =>	x"00000101",
		264 =>	x"01010101",
		265 =>	x"01000101",
		266 =>	x"01000000",
		267 =>	x"00020101",
		268 =>	x"01030101",
		269 =>	x"01000101",
		270 =>	x"01010100",
		271 =>	x"01010202",
		272 =>	x"03030301",
		273 =>	x"01010003",
		274 =>	x"01010101",
		275 =>	x"01010103",
		276 =>	x"02030301",
		277 =>	x"01010003",
		278 =>	x"03030101",
		279 =>	x"01010101",
		280 =>	x"03030301",
		281 =>	x"01010003",
		282 =>	x"03030000",
		283 =>	x"00010103",
		284 =>	x"03030101",
		285 =>	x"03000103",
		286 =>	x"03030000",
		287 =>	x"00010101",
		288 =>	x"01010101",
		289 =>	x"01030301",
		290 =>	x"01030000",
		291 =>	x"00000101",
		292 =>	x"01010101",
		293 =>	x"00010303",
		294 =>	x"01010000",
		295 =>	x"00000000",
		296 =>	x"01000000",
		297 =>	x"00000101",
		298 =>	x"01010202",
		299 =>	x"00000002",
		300 =>	x"00010003",
		301 =>	x"03030303",
		302 =>	x"01020100",
		303 =>	x"00000000",
		304 =>	x"01010101",
		305 =>	x"03030300",
		306 =>	x"00000200",
		307 =>	x"00000000",
		308 =>	x"00000101",
		309 =>	x"01010000",
		310 =>	x"00000000",
		311 =>	x"00000000",
		312 =>	x"00000001",
		313 =>	x"01010100",
		314 =>	x"00000000",
		315 =>	x"00000000",
		316 =>	x"00000000",
		317 =>	x"00010000",
		318 =>	x"00000000",
		319 =>	x"00000000", -- IMG_16x16_avion2_11
		320 =>	x"01010100",
		321 =>	x"00000000",
		322 =>	x"00000000",
		323 =>	x"00000002",
		324 =>	x"01010101",
		325 =>	x"01000000",
		326 =>	x"00000000",
		327 =>	x"00010101",
		328 =>	x"02010101",
		329 =>	x"01010000",
		330 =>	x"00000000",
		331 =>	x"00010101",
		332 =>	x"02030103",
		333 =>	x"01010002",
		334 =>	x"00000000",
		335 =>	x"00010101",
		336 =>	x"03020303",
		337 =>	x"01010100",
		338 =>	x"01000000",
		339 =>	x"01010103",
		340 =>	x"03030303",
		341 =>	x"01010001",
		342 =>	x"01000000",
		343 =>	x"00010101",
		344 =>	x"03030301",
		345 =>	x"01010000",
		346 =>	x"01010000",
		347 =>	x"00000101",
		348 =>	x"01010101",
		349 =>	x"01010003",
		350 =>	x"01010100",
		351 =>	x"00000101",
		352 =>	x"01010103",
		353 =>	x"01000003",
		354 =>	x"03010100",
		355 =>	x"00020000",
		356 =>	x"01010100",
		357 =>	x"03010003",
		358 =>	x"03010101",
		359 =>	x"00010101",
		360 =>	x"00000001",
		361 =>	x"03030103",
		362 =>	x"03000100",
		363 =>	x"00000101",
		364 =>	x"03030303",
		365 =>	x"01030103",
		366 =>	x"00000000",
		367 =>	x"00000101",
		368 =>	x"01030303",
		369 =>	x"01010101",
		370 =>	x"00000000",
		371 =>	x"00000001",
		372 =>	x"01030303",
		373 =>	x"03010102",
		374 =>	x"00000000",
		375 =>	x"00000001",
		376 =>	x"01010000",
		377 =>	x"00000201",
		378 =>	x"02000000",
		379 =>	x"00000000",
		380 =>	x"01010000",
		381 =>	x"00000200",
		382 =>	x"00000000",
		383 =>	x"00000000", -- IMG_16x16_avion2_12
		384 =>	x"00000101",
		385 =>	x"02010100",
		386 =>	x"00000000",
		387 =>	x"00000000",
		388 =>	x"00010101",
		389 =>	x"02010101",
		390 =>	x"00000000",
		391 =>	x"00000000",
		392 =>	x"01010101",
		393 =>	x"02010101",
		394 =>	x"01000000",
		395 =>	x"00000000",
		396 =>	x"01010103",
		397 =>	x"03030101",
		398 =>	x"01000000",
		399 =>	x"00000000",
		400 =>	x"01010303",
		401 =>	x"02030301",
		402 =>	x"01000000",
		403 =>	x"00000000",
		404 =>	x"01010103",
		405 =>	x"03030101",
		406 =>	x"01000000",
		407 =>	x"00000200",
		408 =>	x"01010101",
		409 =>	x"03010101",
		410 =>	x"01000200",
		411 =>	x"00000101",
		412 =>	x"00010101",
		413 =>	x"01010101",
		414 =>	x"00010100",
		415 =>	x"00000101",
		416 =>	x"00000101",
		417 =>	x"03010100",
		418 =>	x"00010100",
		419 =>	x"00000101",
		420 =>	x"03000000",
		421 =>	x"03000000",
		422 =>	x"03010100",
		423 =>	x"00000101",
		424 =>	x"03030001",
		425 =>	x"03010003",
		426 =>	x"03010100",
		427 =>	x"00000101",
		428 =>	x"03030301",
		429 =>	x"03010303",
		430 =>	x"03010100",
		431 =>	x"00000101",
		432 =>	x"00030301",
		433 =>	x"01010303",
		434 =>	x"00010100",
		435 =>	x"00000101",
		436 =>	x"00000301",
		437 =>	x"01010300",
		438 =>	x"00010100",
		439 =>	x"00000000",
		440 =>	x"00000002",
		441 =>	x"01020000",
		442 =>	x"00000000",
		443 =>	x"00000000",
		444 =>	x"00000002",
		445 =>	x"01020000",
		446 =>	x"00000000",
		447 =>	x"00000000", -- IMG_16x16_avion2_9
		448 =>	x"00000000",
		449 =>	x"00000000",
		450 =>	x"00000000",
		451 =>	x"00000000",
		452 =>	x"00000201",
		453 =>	x"01010101",
		454 =>	x"01010000",
		455 =>	x"00000000",
		456 =>	x"00000001",
		457 =>	x"01010101",
		458 =>	x"01010000",
		459 =>	x"00000101",
		460 =>	x"01010100",
		461 =>	x"00030303",
		462 =>	x"00000000",
		463 =>	x"00010101",
		464 =>	x"01010101",
		465 =>	x"00000303",
		466 =>	x"03000000",
		467 =>	x"01010101",
		468 =>	x"03010101",
		469 =>	x"01000003",
		470 =>	x"03030000",
		471 =>	x"01010103",
		472 =>	x"03030101",
		473 =>	x"01000101",
		474 =>	x"01010202",
		475 =>	x"02020203",
		476 =>	x"02030301",
		477 =>	x"03030303",
		478 =>	x"01010101",
		479 =>	x"01010103",
		480 =>	x"03030101",
		481 =>	x"01000101",
		482 =>	x"01010202",
		483 =>	x"01010101",
		484 =>	x"03010101",
		485 =>	x"01000003",
		486 =>	x"03030000",
		487 =>	x"00010101",
		488 =>	x"01010101",
		489 =>	x"00000303",
		490 =>	x"03000000",
		491 =>	x"00000101",
		492 =>	x"01010100",
		493 =>	x"00030303",
		494 =>	x"00000000",
		495 =>	x"00000000",
		496 =>	x"00000001",
		497 =>	x"01010101",
		498 =>	x"01010000",
		499 =>	x"00000000",
		500 =>	x"00000201",
		501 =>	x"01010101",
		502 =>	x"01010000",
		503 =>	x"00000000",
		504 =>	x"00000000",
		505 =>	x"00000000",
		506 =>	x"00000000",
		507 =>	x"00000000",
		508 =>	x"00000000",
		509 =>	x"00000000",
		510 =>	x"00000000",
		511 =>	x"00000000", -- IMG_16x16_avion2_pola10
		512 =>	x"00000000",
		513 =>	x"00000000",
		514 =>	x"00000000",
		515 =>	x"00000000",
		516 =>	x"00000000",
		517 =>	x"02010100",
		518 =>	x"00000000",
		519 =>	x"00000101",
		520 =>	x"01010100",
		521 =>	x"01010101",
		522 =>	x"01010100",
		523 =>	x"00010101",
		524 =>	x"01010101",
		525 =>	x"00000301",
		526 =>	x"01010100",
		527 =>	x"00010101",
		528 =>	x"03030101",
		529 =>	x"01000003",
		530 =>	x"03000000",
		531 =>	x"02020103",
		532 =>	x"03030101",
		533 =>	x"01000003",
		534 =>	x"03000000",
		535 =>	x"01010203",
		536 =>	x"02030301",
		537 =>	x"01000103",
		538 =>	x"03030000",
		539 =>	x"01010103",
		540 =>	x"03030301",
		541 =>	x"03030101",
		542 =>	x"01010000",
		543 =>	x"01010101",
		544 =>	x"03010101",
		545 =>	x"01000303",
		546 =>	x"01010202",
		547 =>	x"00010101",
		548 =>	x"01010101",
		549 =>	x"00000101",
		550 =>	x"01010101",
		551 =>	x"00000101",
		552 =>	x"01010100",
		553 =>	x"00030303",
		554 =>	x"03000202",
		555 =>	x"00000000",
		556 =>	x"00000000",
		557 =>	x"03030303",
		558 =>	x"00000000",
		559 =>	x"00000000",
		560 =>	x"00000101",
		561 =>	x"01030000",
		562 =>	x"00000000",
		563 =>	x"00000000",
		564 =>	x"00020101",
		565 =>	x"01010101",
		566 =>	x"01000000",
		567 =>	x"00000000",
		568 =>	x"00000000",
		569 =>	x"00010101",
		570 =>	x"01000000",
		571 =>	x"00000000",
		572 =>	x"00000000",
		573 =>	x"00000000",
		574 =>	x"00000000",
		575 =>	x"00000101", -- IMG_16x16_avion2_pola11
		576 =>	x"01010100",
		577 =>	x"00000000",
		578 =>	x"00000000",
		579 =>	x"00020101",
		580 =>	x"01010101",
		581 =>	x"00000200",
		582 =>	x"00000000",
		583 =>	x"01010201",
		584 =>	x"01010101",
		585 =>	x"01000101",
		586 =>	x"00000000",
		587 =>	x"01010103",
		588 =>	x"03030301",
		589 =>	x"01000101",
		590 =>	x"01000000",
		591 =>	x"01010103",
		592 =>	x"02030301",
		593 =>	x"01000001",
		594 =>	x"01010000",
		595 =>	x"01010103",
		596 =>	x"03030101",
		597 =>	x"01000303",
		598 =>	x"01010100",
		599 =>	x"01010103",
		600 =>	x"03010301",
		601 =>	x"01000003",
		602 =>	x"03010101",
		603 =>	x"00010101",
		604 =>	x"01010103",
		605 =>	x"00000003",
		606 =>	x"03000101",
		607 =>	x"00000101",
		608 =>	x"01010100",
		609 =>	x"03010103",
		610 =>	x"03000000",
		611 =>	x"00000000",
		612 =>	x"00000000",
		613 =>	x"01030101",
		614 =>	x"03000000",
		615 =>	x"00020101",
		616 =>	x"00030000",
		617 =>	x"01010101",
		618 =>	x"00000000",
		619 =>	x"00000101",
		620 =>	x"01030303",
		621 =>	x"03010101",
		622 =>	x"02000000",
		623 =>	x"00000001",
		624 =>	x"01010303",
		625 =>	x"03030002",
		626 =>	x"01020000",
		627 =>	x"00000000",
		628 =>	x"01010100",
		629 =>	x"00000000",
		630 =>	x"02010000",
		631 =>	x"00000000",
		632 =>	x"00010101",
		633 =>	x"00000000",
		634 =>	x"00000000",
		635 =>	x"00000000",
		636 =>	x"00000101",
		637 =>	x"00000000",
		638 =>	x"00000000",
		639 =>	x"00000000", -- IMG_16x16_avion2_pola12
		640 =>	x"00020101",
		641 =>	x"01000000",
		642 =>	x"00000000",
		643 =>	x"00000001",
		644 =>	x"01020101",
		645 =>	x"01010000",
		646 =>	x"00000000",
		647 =>	x"00000101",
		648 =>	x"01010201",
		649 =>	x"01010100",
		650 =>	x"00000000",
		651 =>	x"00000101",
		652 =>	x"01030303",
		653 =>	x"01010100",
		654 =>	x"00000000",
		655 =>	x"00000101",
		656 =>	x"03030203",
		657 =>	x"03010100",
		658 =>	x"00000000",
		659 =>	x"00000101",
		660 =>	x"03030303",
		661 =>	x"01010100",
		662 =>	x"00020000",
		663 =>	x"00000101",
		664 =>	x"01010303",
		665 =>	x"01010100",
		666 =>	x"01010000",
		667 =>	x"00000001",
		668 =>	x"01010101",
		669 =>	x"01010000",
		670 =>	x"01010000",
		671 =>	x"00020100",
		672 =>	x"01010103",
		673 =>	x"01000003",
		674 =>	x"01010000",
		675 =>	x"00010100",
		676 =>	x"00000003",
		677 =>	x"00000303",
		678 =>	x"03010100",
		679 =>	x"00010103",
		680 =>	x"00000101",
		681 =>	x"03010303",
		682 =>	x"00010100",
		683 =>	x"00000101",
		684 =>	x"03030301",
		685 =>	x"03010303",
		686 =>	x"00010100",
		687 =>	x"00000101",
		688 =>	x"03030301",
		689 =>	x"01010300",
		690 =>	x"00010100",
		691 =>	x"00000101",
		692 =>	x"00000301",
		693 =>	x"01010000",
		694 =>	x"00000000",
		695 =>	x"00000101",
		696 =>	x"00000000",
		697 =>	x"02010200",
		698 =>	x"00000000",
		699 =>	x"00000000",
		700 =>	x"00000000",
		701 =>	x"02010200",
		702 =>	x"00000000",
		703 =>	x"00000000", -- IMG_16x16_avion_10
		704 =>	x"00000000",
		705 =>	x"00000000",
		706 =>	x"00000000",
		707 =>	x"00000000",
		708 =>	x"00000000",
		709 =>	x"00000000",
		710 =>	x"00000000",
		711 =>	x"00000000",
		712 =>	x"00000000",
		713 =>	x"00000004",
		714 =>	x"00000000",
		715 =>	x"00030300",
		716 =>	x"00000004",
		717 =>	x"00000000",
		718 =>	x"04000000",
		719 =>	x"00000303",
		720 =>	x"03030001",
		721 =>	x"03000003",
		722 =>	x"03030300",
		723 =>	x"00000003",
		724 =>	x"03030303",
		725 =>	x"03030303",
		726 =>	x"03030303",
		727 =>	x"00000000",
		728 =>	x"03030304",
		729 =>	x"04030303",
		730 =>	x"00000000",
		731 =>	x"00000000",
		732 =>	x"03030304",
		733 =>	x"03030304",
		734 =>	x"04000000",
		735 =>	x"00000000",
		736 =>	x"00030303",
		737 =>	x"03030303",
		738 =>	x"04000000",
		739 =>	x"00000000",
		740 =>	x"04010303",
		741 =>	x"03030303",
		742 =>	x"00000000",
		743 =>	x"00000000",
		744 =>	x"00030303",
		745 =>	x"03040303",
		746 =>	x"03000000",
		747 =>	x"00000000",
		748 =>	x"00000303",
		749 =>	x"03040400",
		750 =>	x"00000000",
		751 =>	x"00000000",
		752 =>	x"00040003",
		753 =>	x"03000000",
		754 =>	x"00000000",
		755 =>	x"00000000",
		756 =>	x"00000403",
		757 =>	x"03000000",
		758 =>	x"00000000",
		759 =>	x"00000000",
		760 =>	x"00000003",
		761 =>	x"03000000",
		762 =>	x"00000000",
		763 =>	x"00000000",
		764 =>	x"00000000",
		765 =>	x"03030000",
		766 =>	x"00000000",
		767 =>	x"00000000", -- IMG_16x16_avion_11
		768 =>	x"00000000",
		769 =>	x"00000000",
		770 =>	x"00000000",
		771 =>	x"00000003",
		772 =>	x"00000000",
		773 =>	x"00000000",
		774 =>	x"00000000",
		775 =>	x"00000003",
		776 =>	x"03000000",
		777 =>	x"00000000",
		778 =>	x"00000000",
		779 =>	x"00000000",
		780 =>	x"03030000",
		781 =>	x"00000000",
		782 =>	x"00000000",
		783 =>	x"00000000",
		784 =>	x"03030303",
		785 =>	x"00040000",
		786 =>	x"00000000",
		787 =>	x"00000000",
		788 =>	x"03030303",
		789 =>	x"03010300",
		790 =>	x"04000000",
		791 =>	x"00000000",
		792 =>	x"00030303",
		793 =>	x"03030303",
		794 =>	x"00040000",
		795 =>	x"00000004",
		796 =>	x"01030404",
		797 =>	x"03030303",
		798 =>	x"03030300",
		799 =>	x"00000000",
		800 =>	x"03030403",
		801 =>	x"03030303",
		802 =>	x"03030303",
		803 =>	x"00000000",
		804 =>	x"00030303",
		805 =>	x"03030404",
		806 =>	x"00000003",
		807 =>	x"00000000",
		808 =>	x"00030303",
		809 =>	x"03030304",
		810 =>	x"00000000",
		811 =>	x"00000400",
		812 =>	x"03030304",
		813 =>	x"03030300",
		814 =>	x"00000000",
		815 =>	x"00000004",
		816 =>	x"03030004",
		817 =>	x"04000300",
		818 =>	x"00000000",
		819 =>	x"00000000",
		820 =>	x"03030000",
		821 =>	x"00000000",
		822 =>	x"00000000",
		823 =>	x"00000000",
		824 =>	x"03030000",
		825 =>	x"00000000",
		826 =>	x"00000000",
		827 =>	x"00000000",
		828 =>	x"00030000",
		829 =>	x"00000000",
		830 =>	x"00000000",
		831 =>	x"00000000", -- IMG_16x16_avion_12
		832 =>	x"00000000",
		833 =>	x"03000000",
		834 =>	x"00000000",
		835 =>	x"00000000",
		836 =>	x"00000000",
		837 =>	x"03000000",
		838 =>	x"00000000",
		839 =>	x"00000000",
		840 =>	x"00000000",
		841 =>	x"03000000",
		842 =>	x"00000000",
		843 =>	x"00000000",
		844 =>	x"00000003",
		845 =>	x"03030000",
		846 =>	x"00000000",
		847 =>	x"00000000",
		848 =>	x"00000003",
		849 =>	x"03030000",
		850 =>	x"00000000",
		851 =>	x"00000000",
		852 =>	x"04000003",
		853 =>	x"03030000",
		854 =>	x"04000000",
		855 =>	x"00000000",
		856 =>	x"04000003",
		857 =>	x"03030000",
		858 =>	x"04000000",
		859 =>	x"00000000",
		860 =>	x"03000303",
		861 =>	x"03030300",
		862 =>	x"03000000",
		863 =>	x"00040000",
		864 =>	x"03010303",
		865 =>	x"04030301",
		866 =>	x"03000004",
		867 =>	x"00040000",
		868 =>	x"01030304",
		869 =>	x"04040303",
		870 =>	x"01000004",
		871 =>	x"00030000",
		872 =>	x"03030304",
		873 =>	x"03040303",
		874 =>	x"03000003",
		875 =>	x"00030003",
		876 =>	x"03030303",
		877 =>	x"03030303",
		878 =>	x"03030003",
		879 =>	x"00030303",
		880 =>	x"03030403",
		881 =>	x"03030403",
		882 =>	x"03030303",
		883 =>	x"00030303",
		884 =>	x"00040403",
		885 =>	x"03030404",
		886 =>	x"00030303",
		887 =>	x"00030300",
		888 =>	x"00040400",
		889 =>	x"03000404",
		890 =>	x"00000303",
		891 =>	x"00030000",
		892 =>	x"00000000",
		893 =>	x"03000000",
		894 =>	x"00000003",
		895 =>	x"00000000", -- IMG_16x16_avion_9
		896 =>	x"00000000",
		897 =>	x"00000000",
		898 =>	x"00000000",
		899 =>	x"00000000",
		900 =>	x"00000000",
		901 =>	x"04040303",
		902 =>	x"03030303",
		903 =>	x"00000000",
		904 =>	x"00000000",
		905 =>	x"00000000",
		906 =>	x"03030300",
		907 =>	x"00000000",
		908 =>	x"00000000",
		909 =>	x"00000003",
		910 =>	x"03030000",
		911 =>	x"00000000",
		912 =>	x"00040403",
		913 =>	x"03010303",
		914 =>	x"03000000",
		915 =>	x"00000000",
		916 =>	x"00000000",
		917 =>	x"01030303",
		918 =>	x"03040400",
		919 =>	x"00000000",
		920 =>	x"00000003",
		921 =>	x"03030303",
		922 =>	x"04040400",
		923 =>	x"00000003",
		924 =>	x"03030303",
		925 =>	x"03040403",
		926 =>	x"03030000",
		927 =>	x"03030303",
		928 =>	x"03030303",
		929 =>	x"04040303",
		930 =>	x"03030303",
		931 =>	x"00000003",
		932 =>	x"03030303",
		933 =>	x"03040403",
		934 =>	x"03030000",
		935 =>	x"00000000",
		936 =>	x"00000003",
		937 =>	x"03030303",
		938 =>	x"04040400",
		939 =>	x"00000000",
		940 =>	x"00000000",
		941 =>	x"01030303",
		942 =>	x"03040400",
		943 =>	x"00000000",
		944 =>	x"00040403",
		945 =>	x"03010303",
		946 =>	x"03000000",
		947 =>	x"00000000",
		948 =>	x"00000000",
		949 =>	x"00000003",
		950 =>	x"03030000",
		951 =>	x"00000000",
		952 =>	x"00000000",
		953 =>	x"00000000",
		954 =>	x"03030300",
		955 =>	x"00000000",
		956 =>	x"00000000",
		957 =>	x"04040303",
		958 =>	x"03030303",
		959 =>	x"00000000", -- IMG_16x16_avion_pola10
		960 =>	x"00000000",
		961 =>	x"00000000",
		962 =>	x"00000000",
		963 =>	x"00000000",
		964 =>	x"00000000",
		965 =>	x"00000000",
		966 =>	x"00000000",
		967 =>	x"00000000",
		968 =>	x"00000000",
		969 =>	x"00000403",
		970 =>	x"03030000",
		971 =>	x"00000000",
		972 =>	x"00000000",
		973 =>	x"00000000",
		974 =>	x"03030303",
		975 =>	x"00000000",
		976 =>	x"00000403",
		977 =>	x"03010003",
		978 =>	x"03030000",
		979 =>	x"00000003",
		980 =>	x"03000000",
		981 =>	x"01030303",
		982 =>	x"00000000",
		983 =>	x"03030303",
		984 =>	x"03030303",
		985 =>	x"03030303",
		986 =>	x"04040000",
		987 =>	x"00000003",
		988 =>	x"03030304",
		989 =>	x"04040304",
		990 =>	x"04040000",
		991 =>	x"00000000",
		992 =>	x"00030303",
		993 =>	x"04030303",
		994 =>	x"03000000",
		995 =>	x"00000000",
		996 =>	x"00000303",
		997 =>	x"03030303",
		998 =>	x"03030000",
		999 =>	x"00000000",
		1000 =>	x"04030303",
		1001 =>	x"03030404",
		1002 =>	x"04000000",
		1003 =>	x"00000000",
		1004 =>	x"00000001",
		1005 =>	x"03030304",
		1006 =>	x"04000000",
		1007 =>	x"00000000",
		1008 =>	x"00000000",
		1009 =>	x"00030300",
		1010 =>	x"00000000",
		1011 =>	x"00000000",
		1012 =>	x"00000004",
		1013 =>	x"03030300",
		1014 =>	x"00000000",
		1015 =>	x"00000000",
		1016 =>	x"00000000",
		1017 =>	x"00030303",
		1018 =>	x"00000000",
		1019 =>	x"00000000",
		1020 =>	x"00000000",
		1021 =>	x"00000003",
		1022 =>	x"03000000",
		1023 =>	x"00000000", -- IMG_16x16_avion_pola11
		1024 =>	x"00000000",
		1025 =>	x"00000000",
		1026 =>	x"00000000",
		1027 =>	x"00000000",
		1028 =>	x"00000000",
		1029 =>	x"00000000",
		1030 =>	x"00000000",
		1031 =>	x"00030000",
		1032 =>	x"00000000",
		1033 =>	x"00000000",
		1034 =>	x"00000000",
		1035 =>	x"00000300",
		1036 =>	x"00000004",
		1037 =>	x"00000400",
		1038 =>	x"00000000",
		1039 =>	x"00000003",
		1040 =>	x"03000000",
		1041 =>	x"03000004",
		1042 =>	x"00000000",
		1043 =>	x"00000003",
		1044 =>	x"03030000",
		1045 =>	x"01030000",
		1046 =>	x"03000000",
		1047 =>	x"00000000",
		1048 =>	x"03030303",
		1049 =>	x"03030303",
		1050 =>	x"03030000",
		1051 =>	x"00000000",
		1052 =>	x"00030404",
		1053 =>	x"03030303",
		1054 =>	x"03030300",
		1055 =>	x"00000400",
		1056 =>	x"00030403",
		1057 =>	x"03030304",
		1058 =>	x"00000000",
		1059 =>	x"00000003",
		1060 =>	x"01030303",
		1061 =>	x"03030404",
		1062 =>	x"00000000",
		1063 =>	x"00000000",
		1064 =>	x"03030303",
		1065 =>	x"03030000",
		1066 =>	x"00000000",
		1067 =>	x"00000400",
		1068 =>	x"00030303",
		1069 =>	x"04000300",
		1070 =>	x"00000000",
		1071 =>	x"00000004",
		1072 =>	x"00030304",
		1073 =>	x"04000003",
		1074 =>	x"00000000",
		1075 =>	x"00000000",
		1076 =>	x"03030300",
		1077 =>	x"00000000",
		1078 =>	x"00000000",
		1079 =>	x"00000000",
		1080 =>	x"00030300",
		1081 =>	x"00000000",
		1082 =>	x"00000000",
		1083 =>	x"00000000",
		1084 =>	x"00000300",
		1085 =>	x"00000000",
		1086 =>	x"00000000",
		1087 =>	x"00000000", -- IMG_16x16_avion_pola12
		1088 =>	x"00000300",
		1089 =>	x"00000000",
		1090 =>	x"00000000",
		1091 =>	x"00000000",
		1092 =>	x"00000300",
		1093 =>	x"00000000",
		1094 =>	x"00000000",
		1095 =>	x"00000000",
		1096 =>	x"00000300",
		1097 =>	x"00000000",
		1098 =>	x"00000000",
		1099 =>	x"00000000",
		1100 =>	x"00030303",
		1101 =>	x"00000000",
		1102 =>	x"00000000",
		1103 =>	x"00000000",
		1104 =>	x"00030303",
		1105 =>	x"00000400",
		1106 =>	x"00000000",
		1107 =>	x"00000000",
		1108 =>	x"00000303",
		1109 =>	x"03000300",
		1110 =>	x"00000000",
		1111 =>	x"00000000",
		1112 =>	x"04000303",
		1113 =>	x"03030300",
		1114 =>	x"00000000",
		1115 =>	x"00000000",
		1116 =>	x"03000304",
		1117 =>	x"03030301",
		1118 =>	x"00040000",
		1119 =>	x"00000000",
		1120 =>	x"03010304",
		1121 =>	x"04030303",
		1122 =>	x"00030000",
		1123 =>	x"00000000",
		1124 =>	x"01030304",
		1125 =>	x"03030303",
		1126 =>	x"03030300",
		1127 =>	x"00000400",
		1128 =>	x"00030303",
		1129 =>	x"03030403",
		1130 =>	x"03030300",
		1131 =>	x"00000300",
		1132 =>	x"03030304",
		1133 =>	x"03030404",
		1134 =>	x"00000303",
		1135 =>	x"00000303",
		1136 =>	x"03000404",
		1137 =>	x"03030404",
		1138 =>	x"00000003",
		1139 =>	x"00000303",
		1140 =>	x"03000404",
		1141 =>	x"00030000",
		1142 =>	x"00000000",
		1143 =>	x"00000003",
		1144 =>	x"00000000",
		1145 =>	x"00000000",
		1146 =>	x"00000000",
		1147 =>	x"00000003",
		1148 =>	x"00000000",
		1149 =>	x"00000000",
		1150 =>	x"00000000",
		1151 =>	x"00000000", -- IMG_16x16_brod_10
		1152 =>	x"00000000",
		1153 =>	x"00000000",
		1154 =>	x"00000000",
		1155 =>	x"00000000",
		1156 =>	x"00000000",
		1157 =>	x"00000000",
		1158 =>	x"00000000",
		1159 =>	x"00000000",
		1160 =>	x"00000000",
		1161 =>	x"00000003",
		1162 =>	x"00000000",
		1163 =>	x"00020200",
		1164 =>	x"00000003",
		1165 =>	x"00000000",
		1166 =>	x"03000000",
		1167 =>	x"00000202",
		1168 =>	x"02020001",
		1169 =>	x"02000002",
		1170 =>	x"02020200",
		1171 =>	x"00000002",
		1172 =>	x"02020202",
		1173 =>	x"02020202",
		1174 =>	x"02020202",
		1175 =>	x"00000000",
		1176 =>	x"02020203",
		1177 =>	x"03020202",
		1178 =>	x"00000000",
		1179 =>	x"00000000",
		1180 =>	x"02020203",
		1181 =>	x"02020203",
		1182 =>	x"03000000",
		1183 =>	x"00000000",
		1184 =>	x"00020202",
		1185 =>	x"02020202",
		1186 =>	x"03000000",
		1187 =>	x"00000000",
		1188 =>	x"03010202",
		1189 =>	x"02020202",
		1190 =>	x"00000000",
		1191 =>	x"00000000",
		1192 =>	x"00020202",
		1193 =>	x"02030202",
		1194 =>	x"02000000",
		1195 =>	x"00000000",
		1196 =>	x"00000202",
		1197 =>	x"02030300",
		1198 =>	x"00000000",
		1199 =>	x"00000000",
		1200 =>	x"00030002",
		1201 =>	x"02000000",
		1202 =>	x"00000000",
		1203 =>	x"00000000",
		1204 =>	x"00000302",
		1205 =>	x"02000000",
		1206 =>	x"00000000",
		1207 =>	x"00000000",
		1208 =>	x"00000002",
		1209 =>	x"02000000",
		1210 =>	x"00000000",
		1211 =>	x"00000000",
		1212 =>	x"00000000",
		1213 =>	x"02020000",
		1214 =>	x"00000000",
		1215 =>	x"00000000", -- IMG_16x16_brod_11
		1216 =>	x"00000000",
		1217 =>	x"00000000",
		1218 =>	x"00000000",
		1219 =>	x"00000200",
		1220 =>	x"00000000",
		1221 =>	x"00000000",
		1222 =>	x"00000000",
		1223 =>	x"00000202",
		1224 =>	x"00000000",
		1225 =>	x"00000000",
		1226 =>	x"00000000",
		1227 =>	x"00000002",
		1228 =>	x"02000000",
		1229 =>	x"00000000",
		1230 =>	x"00000000",
		1231 =>	x"00000002",
		1232 =>	x"02020200",
		1233 =>	x"03000000",
		1234 =>	x"00000000",
		1235 =>	x"00000002",
		1236 =>	x"02020202",
		1237 =>	x"01020003",
		1238 =>	x"00000000",
		1239 =>	x"00000000",
		1240 =>	x"02020202",
		1241 =>	x"02020200",
		1242 =>	x"03000000",
		1243 =>	x"00000301",
		1244 =>	x"02030302",
		1245 =>	x"02020202",
		1246 =>	x"02020000",
		1247 =>	x"00000002",
		1248 =>	x"02030202",
		1249 =>	x"02020202",
		1250 =>	x"02020200",
		1251 =>	x"00000000",
		1252 =>	x"02020202",
		1253 =>	x"02030300",
		1254 =>	x"00000200",
		1255 =>	x"00000000",
		1256 =>	x"02020202",
		1257 =>	x"02020300",
		1258 =>	x"00000000",
		1259 =>	x"00030002",
		1260 =>	x"02020302",
		1261 =>	x"02020000",
		1262 =>	x"00000000",
		1263 =>	x"00000302",
		1264 =>	x"02000303",
		1265 =>	x"00020000",
		1266 =>	x"00000000",
		1267 =>	x"00000002",
		1268 =>	x"02000000",
		1269 =>	x"00000000",
		1270 =>	x"00000000",
		1271 =>	x"00000002",
		1272 =>	x"02000000",
		1273 =>	x"00000000",
		1274 =>	x"00000000",
		1275 =>	x"00000000",
		1276 =>	x"02000000",
		1277 =>	x"00000000",
		1278 =>	x"00000000",
		1279 =>	x"00000000", -- IMG_16x16_brod_12
		1280 =>	x"00000002",
		1281 =>	x"00000000",
		1282 =>	x"00000000",
		1283 =>	x"00000000",
		1284 =>	x"00000002",
		1285 =>	x"00000000",
		1286 =>	x"00000000",
		1287 =>	x"00000000",
		1288 =>	x"00000002",
		1289 =>	x"00000000",
		1290 =>	x"00000000",
		1291 =>	x"00000000",
		1292 =>	x"00000202",
		1293 =>	x"02000000",
		1294 =>	x"00000000",
		1295 =>	x"00000000",
		1296 =>	x"00000202",
		1297 =>	x"02000000",
		1298 =>	x"00000000",
		1299 =>	x"00000003",
		1300 =>	x"00000202",
		1301 =>	x"02000003",
		1302 =>	x"00000000",
		1303 =>	x"00000003",
		1304 =>	x"00000202",
		1305 =>	x"02000003",
		1306 =>	x"00000000",
		1307 =>	x"00000002",
		1308 =>	x"00020202",
		1309 =>	x"02020002",
		1310 =>	x"00000000",
		1311 =>	x"03000002",
		1312 =>	x"01020203",
		1313 =>	x"02020102",
		1314 =>	x"00000300",
		1315 =>	x"03000001",
		1316 =>	x"02020303",
		1317 =>	x"03020201",
		1318 =>	x"00000300",
		1319 =>	x"02000002",
		1320 =>	x"02020302",
		1321 =>	x"03020202",
		1322 =>	x"00000200",
		1323 =>	x"02000202",
		1324 =>	x"02020202",
		1325 =>	x"02020202",
		1326 =>	x"02000200",
		1327 =>	x"02020202",
		1328 =>	x"02030202",
		1329 =>	x"02030202",
		1330 =>	x"02020200",
		1331 =>	x"02020200",
		1332 =>	x"03030202",
		1333 =>	x"02030300",
		1334 =>	x"02020200",
		1335 =>	x"02020000",
		1336 =>	x"03030002",
		1337 =>	x"00030300",
		1338 =>	x"00020200",
		1339 =>	x"02000000",
		1340 =>	x"00000002",
		1341 =>	x"00000000",
		1342 =>	x"00000200",
		1343 =>	x"00000000", -- IMG_16x16_brod_9
		1344 =>	x"00000000",
		1345 =>	x"00000000",
		1346 =>	x"00000000",
		1347 =>	x"00000000",
		1348 =>	x"00000000",
		1349 =>	x"03030202",
		1350 =>	x"02020202",
		1351 =>	x"00000000",
		1352 =>	x"00000000",
		1353 =>	x"00000000",
		1354 =>	x"02020200",
		1355 =>	x"00000000",
		1356 =>	x"00000000",
		1357 =>	x"00000002",
		1358 =>	x"02020000",
		1359 =>	x"00000000",
		1360 =>	x"00030302",
		1361 =>	x"02010202",
		1362 =>	x"02000000",
		1363 =>	x"00000000",
		1364 =>	x"00000000",
		1365 =>	x"01020202",
		1366 =>	x"02030300",
		1367 =>	x"00000000",
		1368 =>	x"00000002",
		1369 =>	x"02020202",
		1370 =>	x"03030300",
		1371 =>	x"00000002",
		1372 =>	x"02020202",
		1373 =>	x"02030302",
		1374 =>	x"02020000",
		1375 =>	x"02020202",
		1376 =>	x"02020202",
		1377 =>	x"03030202",
		1378 =>	x"02020202",
		1379 =>	x"00000002",
		1380 =>	x"02020202",
		1381 =>	x"02030302",
		1382 =>	x"02020000",
		1383 =>	x"00000000",
		1384 =>	x"00000002",
		1385 =>	x"02020202",
		1386 =>	x"03030300",
		1387 =>	x"00000000",
		1388 =>	x"00000000",
		1389 =>	x"01020202",
		1390 =>	x"02030300",
		1391 =>	x"00000000",
		1392 =>	x"00030302",
		1393 =>	x"02010202",
		1394 =>	x"02000000",
		1395 =>	x"00000000",
		1396 =>	x"00000000",
		1397 =>	x"00000002",
		1398 =>	x"02020000",
		1399 =>	x"00000000",
		1400 =>	x"00000000",
		1401 =>	x"00000000",
		1402 =>	x"02020200",
		1403 =>	x"00000000",
		1404 =>	x"00000000",
		1405 =>	x"03030202",
		1406 =>	x"02020202",
		1407 =>	x"00000000", -- IMG_16x16_brod_pola10
		1408 =>	x"00000000",
		1409 =>	x"00000000",
		1410 =>	x"00000000",
		1411 =>	x"00000000",
		1412 =>	x"00000000",
		1413 =>	x"00000000",
		1414 =>	x"00000000",
		1415 =>	x"00000000",
		1416 =>	x"00000000",
		1417 =>	x"00000000",
		1418 =>	x"00000000",
		1419 =>	x"00000000",
		1420 =>	x"00000000",
		1421 =>	x"00000302",
		1422 =>	x"02020000",
		1423 =>	x"00000000",
		1424 =>	x"00000000",
		1425 =>	x"00000000",
		1426 =>	x"02020202",
		1427 =>	x"00000000",
		1428 =>	x"00000302",
		1429 =>	x"02010002",
		1430 =>	x"02020000",
		1431 =>	x"00000002",
		1432 =>	x"02000000",
		1433 =>	x"01020202",
		1434 =>	x"00000000",
		1435 =>	x"02020202",
		1436 =>	x"02020202",
		1437 =>	x"02020202",
		1438 =>	x"03030000",
		1439 =>	x"00000002",
		1440 =>	x"02020203",
		1441 =>	x"03030203",
		1442 =>	x"03030000",
		1443 =>	x"00000000",
		1444 =>	x"00020202",
		1445 =>	x"03020202",
		1446 =>	x"02000000",
		1447 =>	x"00000000",
		1448 =>	x"00000202",
		1449 =>	x"02020202",
		1450 =>	x"02020000",
		1451 =>	x"00000000",
		1452 =>	x"03020202",
		1453 =>	x"02020303",
		1454 =>	x"03000000",
		1455 =>	x"00000000",
		1456 =>	x"00000001",
		1457 =>	x"02020203",
		1458 =>	x"03000000",
		1459 =>	x"00000000",
		1460 =>	x"00000000",
		1461 =>	x"00020200",
		1462 =>	x"00000000",
		1463 =>	x"00000000",
		1464 =>	x"00000003",
		1465 =>	x"02020200",
		1466 =>	x"00000000",
		1467 =>	x"00000000",
		1468 =>	x"00000000",
		1469 =>	x"00020202",
		1470 =>	x"00000000",
		1471 =>	x"00000000", -- IMG_16x16_brod_pola11
		1472 =>	x"00000000",
		1473 =>	x"00000000",
		1474 =>	x"00000000",
		1475 =>	x"00000000",
		1476 =>	x"00000000",
		1477 =>	x"00000000",
		1478 =>	x"00000000",
		1479 =>	x"00020000",
		1480 =>	x"00000000",
		1481 =>	x"00000000",
		1482 =>	x"00000000",
		1483 =>	x"00000200",
		1484 =>	x"00000003",
		1485 =>	x"00000300",
		1486 =>	x"00000000",
		1487 =>	x"00000002",
		1488 =>	x"02000000",
		1489 =>	x"02000003",
		1490 =>	x"00000000",
		1491 =>	x"00000002",
		1492 =>	x"02020000",
		1493 =>	x"01020000",
		1494 =>	x"02000000",
		1495 =>	x"00000000",
		1496 =>	x"02020202",
		1497 =>	x"02020202",
		1498 =>	x"02020000",
		1499 =>	x"00000000",
		1500 =>	x"00020303",
		1501 =>	x"02020202",
		1502 =>	x"02020200",
		1503 =>	x"00000300",
		1504 =>	x"00020302",
		1505 =>	x"02020203",
		1506 =>	x"00000000",
		1507 =>	x"00000002",
		1508 =>	x"01020202",
		1509 =>	x"02020303",
		1510 =>	x"00000000",
		1511 =>	x"00000000",
		1512 =>	x"02020202",
		1513 =>	x"02020000",
		1514 =>	x"00000000",
		1515 =>	x"00000300",
		1516 =>	x"00020202",
		1517 =>	x"03000200",
		1518 =>	x"00000000",
		1519 =>	x"00000003",
		1520 =>	x"00020203",
		1521 =>	x"03000002",
		1522 =>	x"00000000",
		1523 =>	x"00000000",
		1524 =>	x"02020200",
		1525 =>	x"00000000",
		1526 =>	x"00000000",
		1527 =>	x"00000000",
		1528 =>	x"00020200",
		1529 =>	x"00000000",
		1530 =>	x"00000000",
		1531 =>	x"00000000",
		1532 =>	x"00000200",
		1533 =>	x"00000000",
		1534 =>	x"00000000",
		1535 =>	x"00000000", -- IMG_16x16_brod_pola12
		1536 =>	x"00020000",
		1537 =>	x"00000000",
		1538 =>	x"00000000",
		1539 =>	x"00000000",
		1540 =>	x"00020000",
		1541 =>	x"00000000",
		1542 =>	x"00000000",
		1543 =>	x"00000000",
		1544 =>	x"00020000",
		1545 =>	x"00000000",
		1546 =>	x"00000000",
		1547 =>	x"00000000",
		1548 =>	x"02020200",
		1549 =>	x"00000000",
		1550 =>	x"00000000",
		1551 =>	x"00000000",
		1552 =>	x"02020200",
		1553 =>	x"00030000",
		1554 =>	x"00000000",
		1555 =>	x"00000000",
		1556 =>	x"00020202",
		1557 =>	x"00020000",
		1558 =>	x"00000000",
		1559 =>	x"00000003",
		1560 =>	x"00020202",
		1561 =>	x"02020000",
		1562 =>	x"00000000",
		1563 =>	x"00000002",
		1564 =>	x"00020302",
		1565 =>	x"02020100",
		1566 =>	x"03000000",
		1567 =>	x"00000002",
		1568 =>	x"01020303",
		1569 =>	x"02020200",
		1570 =>	x"02000000",
		1571 =>	x"00000001",
		1572 =>	x"02020302",
		1573 =>	x"02020202",
		1574 =>	x"02020000",
		1575 =>	x"00030000",
		1576 =>	x"02020202",
		1577 =>	x"02030202",
		1578 =>	x"02020000",
		1579 =>	x"00020002",
		1580 =>	x"02020302",
		1581 =>	x"02030300",
		1582 =>	x"00020200",
		1583 =>	x"00020202",
		1584 =>	x"00030302",
		1585 =>	x"02030300",
		1586 =>	x"00000200",
		1587 =>	x"00020202",
		1588 =>	x"00030300",
		1589 =>	x"02000000",
		1590 =>	x"00000000",
		1591 =>	x"00000200",
		1592 =>	x"00000000",
		1593 =>	x"00000000",
		1594 =>	x"00000000",
		1595 =>	x"00000200",
		1596 =>	x"00000000",
		1597 =>	x"00000000",
		1598 =>	x"00000000",
		1599 =>	x"00000000", -- IMG_16x16_crno
		1600 =>	x"00000000",
		1601 =>	x"00000000",
		1602 =>	x"00000000",
		1603 =>	x"00000000",
		1604 =>	x"00000000",
		1605 =>	x"00000000",
		1606 =>	x"00000000",
		1607 =>	x"00000000",
		1608 =>	x"00000000",
		1609 =>	x"00000000",
		1610 =>	x"00000000",
		1611 =>	x"00000000",
		1612 =>	x"00000000",
		1613 =>	x"00000000",
		1614 =>	x"00000000",
		1615 =>	x"00000000",
		1616 =>	x"00000000",
		1617 =>	x"00000000",
		1618 =>	x"00000000",
		1619 =>	x"00000000",
		1620 =>	x"00000000",
		1621 =>	x"00000000",
		1622 =>	x"00000000",
		1623 =>	x"00000000",
		1624 =>	x"00000000",
		1625 =>	x"00000000",
		1626 =>	x"00000000",
		1627 =>	x"00000000",
		1628 =>	x"00000000",
		1629 =>	x"00000000",
		1630 =>	x"00000000",
		1631 =>	x"00000000",
		1632 =>	x"00000000",
		1633 =>	x"00000000",
		1634 =>	x"00000000",
		1635 =>	x"00000000",
		1636 =>	x"00000000",
		1637 =>	x"00000000",
		1638 =>	x"00000000",
		1639 =>	x"00000000",
		1640 =>	x"00000000",
		1641 =>	x"00000000",
		1642 =>	x"00000000",
		1643 =>	x"00000000",
		1644 =>	x"00000000",
		1645 =>	x"00000000",
		1646 =>	x"00000000",
		1647 =>	x"00000000",
		1648 =>	x"00000000",
		1649 =>	x"00000000",
		1650 =>	x"00000000",
		1651 =>	x"00000000",
		1652 =>	x"00000000",
		1653 =>	x"00000000",
		1654 =>	x"00000000",
		1655 =>	x"00000000",
		1656 =>	x"00000000",
		1657 =>	x"00000000",
		1658 =>	x"00000000",
		1659 =>	x"00000000",
		1660 =>	x"00000000",
		1661 =>	x"00000000",
		1662 =>	x"00000000",
		1663 =>	x"00000000", -- IMG_16x16_metak_12
		1664 =>	x"00000000",
		1665 =>	x"00000000",
		1666 =>	x"00000000",
		1667 =>	x"00000000",
		1668 =>	x"00000000",
		1669 =>	x"00000000",
		1670 =>	x"00000000",
		1671 =>	x"00000000",
		1672 =>	x"00000000",
		1673 =>	x"00000000",
		1674 =>	x"00000000",
		1675 =>	x"00000000",
		1676 =>	x"00000000",
		1677 =>	x"00000000",
		1678 =>	x"00000000",
		1679 =>	x"00000000",
		1680 =>	x"00000005",
		1681 =>	x"05000000",
		1682 =>	x"00000000",
		1683 =>	x"00000000",
		1684 =>	x"00000005",
		1685 =>	x"05000000",
		1686 =>	x"00000000",
		1687 =>	x"00000000",
		1688 =>	x"00000505",
		1689 =>	x"05050000",
		1690 =>	x"00000000",
		1691 =>	x"00000000",
		1692 =>	x"00000506",
		1693 =>	x"06050000",
		1694 =>	x"00000000",
		1695 =>	x"00000000",
		1696 =>	x"00000006",
		1697 =>	x"06000000",
		1698 =>	x"00000000",
		1699 =>	x"00000000",
		1700 =>	x"00000006",
		1701 =>	x"06000000",
		1702 =>	x"00000000",
		1703 =>	x"00000000",
		1704 =>	x"00000006",
		1705 =>	x"06000000",
		1706 =>	x"00000000",
		1707 =>	x"00000000",
		1708 =>	x"00000006",
		1709 =>	x"06000000",
		1710 =>	x"00000000",
		1711 =>	x"00000000",
		1712 =>	x"00000000",
		1713 =>	x"00000000",
		1714 =>	x"00000000",
		1715 =>	x"00000000",
		1716 =>	x"00000000",
		1717 =>	x"00000000",
		1718 =>	x"00000000",
		1719 =>	x"00000000",
		1720 =>	x"00000000",
		1721 =>	x"00000000",
		1722 =>	x"00000000",
		1723 =>	x"00000000",
		1724 =>	x"00000000",
		1725 =>	x"00000000",
		1726 =>	x"00000000",
		1727 =>	x"00000000", -- IMG_16x16_metak_muva_12
		1728 =>	x"00000000",
		1729 =>	x"00000000",
		1730 =>	x"00000000",
		1731 =>	x"00000000",
		1732 =>	x"00000000",
		1733 =>	x"00000000",
		1734 =>	x"00000000",
		1735 =>	x"00000000",
		1736 =>	x"00000000",
		1737 =>	x"00000000",
		1738 =>	x"00000000",
		1739 =>	x"00000000",
		1740 =>	x"00000000",
		1741 =>	x"00000000",
		1742 =>	x"00000000",
		1743 =>	x"00000000",
		1744 =>	x"00000006",
		1745 =>	x"00000000",
		1746 =>	x"00000000",
		1747 =>	x"00000000",
		1748 =>	x"00000006",
		1749 =>	x"00000000",
		1750 =>	x"00000000",
		1751 =>	x"00000000",
		1752 =>	x"00000606",
		1753 =>	x"06000000",
		1754 =>	x"00000000",
		1755 =>	x"00000000",
		1756 =>	x"00000607",
		1757 =>	x"06000000",
		1758 =>	x"00000000",
		1759 =>	x"00000000",
		1760 =>	x"00000008",
		1761 =>	x"00000000",
		1762 =>	x"00000000",
		1763 =>	x"00000000",
		1764 =>	x"00000008",
		1765 =>	x"00000000",
		1766 =>	x"00000000",
		1767 =>	x"00000000",
		1768 =>	x"00000008",
		1769 =>	x"00000000",
		1770 =>	x"00000000",
		1771 =>	x"00000000",
		1772 =>	x"00000008",
		1773 =>	x"00000000",
		1774 =>	x"00000000",
		1775 =>	x"00000000",
		1776 =>	x"00000000",
		1777 =>	x"00000000",
		1778 =>	x"00000000",
		1779 =>	x"00000000",
		1780 =>	x"00000000",
		1781 =>	x"00000000",
		1782 =>	x"00000000",
		1783 =>	x"00000000",
		1784 =>	x"00000000",
		1785 =>	x"00000000",
		1786 =>	x"00000000",
		1787 =>	x"00000000",
		1788 =>	x"00000000",
		1789 =>	x"00000000",
		1790 =>	x"00000000",
		1791 =>	x"00000000", -- IMG_16x16_muva2_10
		1792 =>	x"00000000",
		1793 =>	x"00000000",
		1794 =>	x"00000000",
		1795 =>	x"00000000",
		1796 =>	x"01000000",
		1797 =>	x"00010000",
		1798 =>	x"00000000",
		1799 =>	x"00000000",
		1800 =>	x"01000000",
		1801 =>	x"01010000",
		1802 =>	x"00000000",
		1803 =>	x"00000109",
		1804 =>	x"09010001",
		1805 =>	x"01010101",
		1806 =>	x"01010000",
		1807 =>	x"00010101",
		1808 =>	x"01010A01",
		1809 =>	x"01010909",
		1810 =>	x"09010100",
		1811 =>	x"00000909",
		1812 =>	x"010A0A0A",
		1813 =>	x"0A010101",
		1814 =>	x"09010101",
		1815 =>	x"00000901",
		1816 =>	x"0A0A0A0A",
		1817 =>	x"09000000",
		1818 =>	x"01010100",
		1819 =>	x"00010100",
		1820 =>	x"0A0A0A0A",
		1821 =>	x"00000000",
		1822 =>	x"00000000",
		1823 =>	x"00000000",
		1824 =>	x"010A0A09",
		1825 =>	x"09000000",
		1826 =>	x"00000000",
		1827 =>	x"00000001",
		1828 =>	x"01010100",
		1829 =>	x"00000000",
		1830 =>	x"00000000",
		1831 =>	x"00000001",
		1832 =>	x"01010100",
		1833 =>	x"00000000",
		1834 =>	x"00000000",
		1835 =>	x"00000001",
		1836 =>	x"01010101",
		1837 =>	x"01000000",
		1838 =>	x"00000000",
		1839 =>	x"00000000",
		1840 =>	x"00010101",
		1841 =>	x"09010100",
		1842 =>	x"00000000",
		1843 =>	x"00000000",
		1844 =>	x"00000109",
		1845 =>	x"09010100",
		1846 =>	x"00000000",
		1847 =>	x"00000000",
		1848 =>	x"00000001",
		1849 =>	x"01010100",
		1850 =>	x"00000000",
		1851 =>	x"00000000",
		1852 =>	x"00000000",
		1853 =>	x"00000000",
		1854 =>	x"00000000",
		1855 =>	x"00000000", -- IMG_16x16_muva2_11
		1856 =>	x"00000000",
		1857 =>	x"00000000",
		1858 =>	x"00000000",
		1859 =>	x"00000000",
		1860 =>	x"01000001",
		1861 =>	x"00000000",
		1862 =>	x"00000000",
		1863 =>	x"00000001",
		1864 =>	x"01090901",
		1865 =>	x"00000000",
		1866 =>	x"00000000",
		1867 =>	x"00000009",
		1868 =>	x"01090100",
		1869 =>	x"00010101",
		1870 =>	x"00000000",
		1871 =>	x"00010109",
		1872 =>	x"01010A0A",
		1873 =>	x"01010101",
		1874 =>	x"00000000",
		1875 =>	x"00000001",
		1876 =>	x"010A0A0A",
		1877 =>	x"0A010101",
		1878 =>	x"01000000",
		1879 =>	x"00000000",
		1880 =>	x"0A0A0A0A",
		1881 =>	x"0A010101",
		1882 =>	x"01010000",
		1883 =>	x"00000001",
		1884 =>	x"010A0A0A",
		1885 =>	x"09000001",
		1886 =>	x"01090100",
		1887 =>	x"00000101",
		1888 =>	x"010A0900",
		1889 =>	x"09000001",
		1890 =>	x"09090100",
		1891 =>	x"00010101",
		1892 =>	x"01010000",
		1893 =>	x"00000000",
		1894 =>	x"01010100",
		1895 =>	x"00000001",
		1896 =>	x"09010000",
		1897 =>	x"00000000",
		1898 =>	x"01010100",
		1899 =>	x"00000001",
		1900 =>	x"09010000",
		1901 =>	x"00000000",
		1902 =>	x"00000000",
		1903 =>	x"00000001",
		1904 =>	x"09090100",
		1905 =>	x"00000000",
		1906 =>	x"00000000",
		1907 =>	x"00000001",
		1908 =>	x"01010100",
		1909 =>	x"00000000",
		1910 =>	x"00000000",
		1911 =>	x"00000000",
		1912 =>	x"01010100",
		1913 =>	x"00000000",
		1914 =>	x"00000000",
		1915 =>	x"00000000",
		1916 =>	x"00010000",
		1917 =>	x"00000000",
		1918 =>	x"00000000",
		1919 =>	x"00000000", -- IMG_16x16_muva2_12_rasireno
		1920 =>	x"00000001",
		1921 =>	x"00010000",
		1922 =>	x"00000000",
		1923 =>	x"00000000",
		1924 =>	x"00000001",
		1925 =>	x"00010000",
		1926 =>	x"00000000",
		1927 =>	x"00000000",
		1928 =>	x"01010909",
		1929 =>	x"01090901",
		1930 =>	x"01000000",
		1931 =>	x"00000000",
		1932 =>	x"00010909",
		1933 =>	x"01090901",
		1934 =>	x"00000000",
		1935 =>	x"00000000",
		1936 =>	x"00000101",
		1937 =>	x"01010100",
		1938 =>	x"00000000",
		1939 =>	x"00000000",
		1940 =>	x"00010A0A",
		1941 =>	x"010A0A01",
		1942 =>	x"00000000",
		1943 =>	x"00000001",
		1944 =>	x"01010A0A",
		1945 =>	x"0A0A0A01",
		1946 =>	x"01010000",
		1947 =>	x"00010101",
		1948 =>	x"01010A0A",
		1949 =>	x"0A0A0A01",
		1950 =>	x"01010101",
		1951 =>	x"00000101",
		1952 =>	x"01010A0A",
		1953 =>	x"0A0A0A01",
		1954 =>	x"01010100",
		1955 =>	x"00000109",
		1956 =>	x"01010009",
		1957 =>	x"00090001",
		1958 =>	x"01090100",
		1959 =>	x"00010109",
		1960 =>	x"01000009",
		1961 =>	x"00090000",
		1962 =>	x"01090101",
		1963 =>	x"00010901",
		1964 =>	x"01000000",
		1965 =>	x"00000000",
		1966 =>	x"01010901",
		1967 =>	x"00010909",
		1968 =>	x"01000000",
		1969 =>	x"00000000",
		1970 =>	x"01090901",
		1971 =>	x"00010909",
		1972 =>	x"01000000",
		1973 =>	x"00000000",
		1974 =>	x"01090901",
		1975 =>	x"00010101",
		1976 =>	x"01000000",
		1977 =>	x"00000000",
		1978 =>	x"01010101",
		1979 =>	x"00000101",
		1980 =>	x"00000000",
		1981 =>	x"00000000",
		1982 =>	x"00010100",
		1983 =>	x"00000000", -- IMG_16x16_muva2_12_skupljeno
		1984 =>	x"00000000",
		1985 =>	x"00000000",
		1986 =>	x"00000000",
		1987 =>	x"00000000",
		1988 =>	x"00000001",
		1989 =>	x"00010000",
		1990 =>	x"00000000",
		1991 =>	x"00000000",
		1992 =>	x"01010909",
		1993 =>	x"01090901",
		1994 =>	x"01000000",
		1995 =>	x"00000000",
		1996 =>	x"00010909",
		1997 =>	x"01090901",
		1998 =>	x"00000000",
		1999 =>	x"00000000",
		2000 =>	x"00000101",
		2001 =>	x"01010100",
		2002 =>	x"00000000",
		2003 =>	x"00000000",
		2004 =>	x"01010A0A",
		2005 =>	x"010A0A01",
		2006 =>	x"01000000",
		2007 =>	x"00000001",
		2008 =>	x"01010A0A",
		2009 =>	x"0A0A0A01",
		2010 =>	x"01010000",
		2011 =>	x"00010101",
		2012 =>	x"01010A0A",
		2013 =>	x"0A0A0A01",
		2014 =>	x"01010101",
		2015 =>	x"00000101",
		2016 =>	x"01000A0A",
		2017 =>	x"0A0A0A00",
		2018 =>	x"01010100",
		2019 =>	x"00000001",
		2020 =>	x"01000009",
		2021 =>	x"00090000",
		2022 =>	x"01010000",
		2023 =>	x"00000001",
		2024 =>	x"01000009",
		2025 =>	x"00090000",
		2026 =>	x"01010000",
		2027 =>	x"00000001",
		2028 =>	x"01010000",
		2029 =>	x"00000001",
		2030 =>	x"01010000",
		2031 =>	x"00000000",
		2032 =>	x"01010000",
		2033 =>	x"00000001",
		2034 =>	x"01000000",
		2035 =>	x"00000000",
		2036 =>	x"00010100",
		2037 =>	x"00000101",
		2038 =>	x"00000000",
		2039 =>	x"00000000",
		2040 =>	x"00000101",
		2041 =>	x"00010100",
		2042 =>	x"00000000",
		2043 =>	x"00000000",
		2044 =>	x"00000001",
		2045 =>	x"00010000",
		2046 =>	x"00000000",
		2047 =>	x"00000000", -- IMG_16x16_muva2_9
		2048 =>	x"00000000",
		2049 =>	x"00000000",
		2050 =>	x"00000000",
		2051 =>	x"00000000",
		2052 =>	x"00000001",
		2053 =>	x"00000101",
		2054 =>	x"01010100",
		2055 =>	x"00000000",
		2056 =>	x"00000001",
		2057 =>	x"01010109",
		2058 =>	x"09090101",
		2059 =>	x"00000000",
		2060 =>	x"00000101",
		2061 =>	x"01090901",
		2062 =>	x"09090101",
		2063 =>	x"00000100",
		2064 =>	x"00000101",
		2065 =>	x"01010101",
		2066 =>	x"01010100",
		2067 =>	x"00000101",
		2068 =>	x"00010101",
		2069 =>	x"01010000",
		2070 =>	x"00000000",
		2071 =>	x"00000909",
		2072 =>	x"010A0A0A",
		2073 =>	x"0A000000",
		2074 =>	x"00000000",
		2075 =>	x"01010909",
		2076 =>	x"010A0A0A",
		2077 =>	x"0A090900",
		2078 =>	x"00000000",
		2079 =>	x"00000101",
		2080 =>	x"01010A0A",
		2081 =>	x"0A000000",
		2082 =>	x"00000000",
		2083 =>	x"01010909",
		2084 =>	x"010A0A0A",
		2085 =>	x"0A090900",
		2086 =>	x"00000000",
		2087 =>	x"00000909",
		2088 =>	x"010A0A0A",
		2089 =>	x"0A000000",
		2090 =>	x"00000000",
		2091 =>	x"00000101",
		2092 =>	x"00010101",
		2093 =>	x"01010000",
		2094 =>	x"00000000",
		2095 =>	x"00000100",
		2096 =>	x"00000101",
		2097 =>	x"01010101",
		2098 =>	x"01010100",
		2099 =>	x"00000000",
		2100 =>	x"00000101",
		2101 =>	x"01090901",
		2102 =>	x"09090101",
		2103 =>	x"00000000",
		2104 =>	x"00000001",
		2105 =>	x"01010109",
		2106 =>	x"09090101",
		2107 =>	x"00000000",
		2108 =>	x"00000001",
		2109 =>	x"00000101",
		2110 =>	x"01010100",
		2111 =>	x"00000000", -- IMG_16x16_muva2_pola10
		2112 =>	x"00000000",
		2113 =>	x"00000000",
		2114 =>	x"00000000",
		2115 =>	x"00000000",
		2116 =>	x"00000000",
		2117 =>	x"00010000",
		2118 =>	x"00000000",
		2119 =>	x"00000001",
		2120 =>	x"00000000",
		2121 =>	x"01010100",
		2122 =>	x"00000000",
		2123 =>	x"00000001",
		2124 =>	x"01000101",
		2125 =>	x"01010101",
		2126 =>	x"01000000",
		2127 =>	x"00000009",
		2128 =>	x"01000101",
		2129 =>	x"01010101",
		2130 =>	x"01000000",
		2131 =>	x"00000109",
		2132 =>	x"09010A0A",
		2133 =>	x"01000000",
		2134 =>	x"01010000",
		2135 =>	x"00000101",
		2136 =>	x"010A0A0A",
		2137 =>	x"0A0A0000",
		2138 =>	x"01010100",
		2139 =>	x"00010909",
		2140 =>	x"01010A0A",
		2141 =>	x"0A090900",
		2142 =>	x"00010100",
		2143 =>	x"00000909",
		2144 =>	x"010A0A0A",
		2145 =>	x"0A000000",
		2146 =>	x"00000101",
		2147 =>	x"00000100",
		2148 =>	x"010A0A0A",
		2149 =>	x"0A090900",
		2150 =>	x"00000000",
		2151 =>	x"00010000",
		2152 =>	x"0101010A",
		2153 =>	x"00000000",
		2154 =>	x"00000100",
		2155 =>	x"00000000",
		2156 =>	x"01010100",
		2157 =>	x"00000100",
		2158 =>	x"01010000",
		2159 =>	x"00000000",
		2160 =>	x"00010101",
		2161 =>	x"01010101",
		2162 =>	x"01000000",
		2163 =>	x"00000000",
		2164 =>	x"00000101",
		2165 =>	x"01010101",
		2166 =>	x"00000000",
		2167 =>	x"00000000",
		2168 =>	x"00010000",
		2169 =>	x"00000000",
		2170 =>	x"00000000",
		2171 =>	x"00000000",
		2172 =>	x"00000000",
		2173 =>	x"00000000",
		2174 =>	x"00000000",
		2175 =>	x"00000000", -- IMG_16x16_muva2_pola11
		2176 =>	x"00000000",
		2177 =>	x"00000000",
		2178 =>	x"00000000",
		2179 =>	x"00000000",
		2180 =>	x"00000001",
		2181 =>	x"00000000",
		2182 =>	x"00000000",
		2183 =>	x"00000000",
		2184 =>	x"00000001",
		2185 =>	x"00000000",
		2186 =>	x"00000000",
		2187 =>	x"00000000",
		2188 =>	x"01090900",
		2189 =>	x"00010100",
		2190 =>	x"01010000",
		2191 =>	x"00000001",
		2192 =>	x"00090901",
		2193 =>	x"01010101",
		2194 =>	x"01000000",
		2195 =>	x"00000009",
		2196 =>	x"0901010A",
		2197 =>	x"0A010101",
		2198 =>	x"01000000",
		2199 =>	x"00000009",
		2200 =>	x"0901010A",
		2201 =>	x"0A0A0001",
		2202 =>	x"01010000",
		2203 =>	x"00010100",
		2204 =>	x"010A0A0A",
		2205 =>	x"0A0A0A00",
		2206 =>	x"01010100",
		2207 =>	x"00000000",
		2208 =>	x"010A0A0A",
		2209 =>	x"0A0A0900",
		2210 =>	x"01010100",
		2211 =>	x"00000001",
		2212 =>	x"01010A0A",
		2213 =>	x"0A000900",
		2214 =>	x"00010100",
		2215 =>	x"00000001",
		2216 =>	x"0101000A",
		2217 =>	x"09090000",
		2218 =>	x"00010100",
		2219 =>	x"00000000",
		2220 =>	x"01010100",
		2221 =>	x"00000000",
		2222 =>	x"00010000",
		2223 =>	x"00000001",
		2224 =>	x"01010101",
		2225 =>	x"01000000",
		2226 =>	x"00010000",
		2227 =>	x"00000001",
		2228 =>	x"00000101",
		2229 =>	x"01010101",
		2230 =>	x"01000000",
		2231 =>	x"00000000",
		2232 =>	x"00000001",
		2233 =>	x"01010100",
		2234 =>	x"00000000",
		2235 =>	x"00000000",
		2236 =>	x"00000000",
		2237 =>	x"00000000",
		2238 =>	x"00000000",
		2239 =>	x"00000000", -- IMG_16x16_muva2_pola12
		2240 =>	x"00000000",
		2241 =>	x"00000000",
		2242 =>	x"00000000",
		2243 =>	x"00000000",
		2244 =>	x"00000001",
		2245 =>	x"00000100",
		2246 =>	x"00000000",
		2247 =>	x"00000000",
		2248 =>	x"00010109",
		2249 =>	x"09010000",
		2250 =>	x"00000000",
		2251 =>	x"00000101",
		2252 =>	x"09090109",
		2253 =>	x"09000000",
		2254 =>	x"00000000",
		2255 =>	x"00000001",
		2256 =>	x"01090101",
		2257 =>	x"01010101",
		2258 =>	x"00000000",
		2259 =>	x"00000000",
		2260 =>	x"00010A01",
		2261 =>	x"0A0A0101",
		2262 =>	x"01000100",
		2263 =>	x"00000001",
		2264 =>	x"010A0A0A",
		2265 =>	x"0A0A0101",
		2266 =>	x"01010000",
		2267 =>	x"00000001",
		2268 =>	x"010A0A0A",
		2269 =>	x"0A0A0A00",
		2270 =>	x"01010000",
		2271 =>	x"00000101",
		2272 =>	x"01010A0A",
		2273 =>	x"0A0A0000",
		2274 =>	x"01010000",
		2275 =>	x"00010101",
		2276 =>	x"01000A09",
		2277 =>	x"00090000",
		2278 =>	x"01010000",
		2279 =>	x"00000101",
		2280 =>	x"01000009",
		2281 =>	x"00090001",
		2282 =>	x"01010000",
		2283 =>	x"00000001",
		2284 =>	x"01000000",
		2285 =>	x"00000000",
		2286 =>	x"01010000",
		2287 =>	x"00000001",
		2288 =>	x"01010100",
		2289 =>	x"00000001",
		2290 =>	x"01000000",
		2291 =>	x"00000000",
		2292 =>	x"00010101",
		2293 =>	x"00000001",
		2294 =>	x"00000000",
		2295 =>	x"00000000",
		2296 =>	x"00000101",
		2297 =>	x"01000100",
		2298 =>	x"00000000",
		2299 =>	x"00000000",
		2300 =>	x"00000000",
		2301 =>	x"01000000",
		2302 =>	x"00000000",
		2303 =>	x"00000000", -- IMG_16x16_muva3_10
		2304 =>	x"00000000",
		2305 =>	x"00000000",
		2306 =>	x"00000000",
		2307 =>	x"00000000",
		2308 =>	x"00000003",
		2309 =>	x"03030000",
		2310 =>	x"00000000",
		2311 =>	x"00000000",
		2312 =>	x"00000303",
		2313 =>	x"03030000",
		2314 =>	x"00000000",
		2315 =>	x"00000000",
		2316 =>	x"00000003",
		2317 =>	x"03030300",
		2318 =>	x"00000000",
		2319 =>	x"00000000",
		2320 =>	x"01000000",
		2321 =>	x"00030303",
		2322 =>	x"03000000",
		2323 =>	x"00000000",
		2324 =>	x"00010302",
		2325 =>	x"03030303",
		2326 =>	x"03000000",
		2327 =>	x"00000001",
		2328 =>	x"00000202",
		2329 =>	x"03030303",
		2330 =>	x"03000000",
		2331 =>	x"00000000",
		2332 =>	x"01030202",
		2333 =>	x"02010303",
		2334 =>	x"03030000",
		2335 =>	x"00000000",
		2336 =>	x"00020202",
		2337 =>	x"01010202",
		2338 =>	x"00000000",
		2339 =>	x"00000303",
		2340 =>	x"00000303",
		2341 =>	x"01020201",
		2342 =>	x"00000000",
		2343 =>	x"00000003",
		2344 =>	x"03000303",
		2345 =>	x"03020101",
		2346 =>	x"01000000",
		2347 =>	x"00000303",
		2348 =>	x"03030303",
		2349 =>	x"03030000",
		2350 =>	x"00000000",
		2351 =>	x"00000003",
		2352 =>	x"03030303",
		2353 =>	x"03030300",
		2354 =>	x"00000000",
		2355 =>	x"00000000",
		2356 =>	x"00000003",
		2357 =>	x"03030000",
		2358 =>	x"00000000",
		2359 =>	x"00000000",
		2360 =>	x"00000003",
		2361 =>	x"00030000",
		2362 =>	x"00000000",
		2363 =>	x"00000000",
		2364 =>	x"00000000",
		2365 =>	x"00000000",
		2366 =>	x"00000000",
		2367 =>	x"00000000", -- IMG_16x16_muva3_11
		2368 =>	x"00000000",
		2369 =>	x"00000000",
		2370 =>	x"00000000",
		2371 =>	x"00000000",
		2372 =>	x"00000000",
		2373 =>	x"00000000",
		2374 =>	x"00000000",
		2375 =>	x"00000000",
		2376 =>	x"00000000",
		2377 =>	x"00030003",
		2378 =>	x"00000000",
		2379 =>	x"00000000",
		2380 =>	x"00000100",
		2381 =>	x"00030303",
		2382 =>	x"03000000",
		2383 =>	x"00000000",
		2384 =>	x"01000001",
		2385 =>	x"00000303",
		2386 =>	x"03000000",
		2387 =>	x"00000000",
		2388 =>	x"00010003",
		2389 =>	x"02000003",
		2390 =>	x"03000000",
		2391 =>	x"00000300",
		2392 =>	x"00030202",
		2393 =>	x"02030303",
		2394 =>	x"03000000",
		2395 =>	x"00030303",
		2396 =>	x"00020202",
		2397 =>	x"02030303",
		2398 =>	x"03030300",
		2399 =>	x"00030303",
		2400 =>	x"00030302",
		2401 =>	x"01010303",
		2402 =>	x"03030000",
		2403 =>	x"00030303",
		2404 =>	x"03030301",
		2405 =>	x"01020203",
		2406 =>	x"03030300",
		2407 =>	x"00000003",
		2408 =>	x"03030303",
		2409 =>	x"02020100",
		2410 =>	x"03000000",
		2411 =>	x"00000000",
		2412 =>	x"03030303",
		2413 =>	x"02010100",
		2414 =>	x"00000000",
		2415 =>	x"00000000",
		2416 =>	x"03030303",
		2417 =>	x"00000100",
		2418 =>	x"00000000",
		2419 =>	x"00000000",
		2420 =>	x"00000003",
		2421 =>	x"00000000",
		2422 =>	x"00000000",
		2423 =>	x"00000000",
		2424 =>	x"00000000",
		2425 =>	x"00000000",
		2426 =>	x"00000000",
		2427 =>	x"00000000",
		2428 =>	x"00000000",
		2429 =>	x"00000000",
		2430 =>	x"00000000",
		2431 =>	x"00000000", -- IMG_16x16_muva3_12_rasireno
		2432 =>	x"00000000",
		2433 =>	x"00000000",
		2434 =>	x"00000000",
		2435 =>	x"00000000",
		2436 =>	x"00000000",
		2437 =>	x"00000000",
		2438 =>	x"00000000",
		2439 =>	x"00000000",
		2440 =>	x"00000000",
		2441 =>	x"00000000",
		2442 =>	x"00000000",
		2443 =>	x"00000000",
		2444 =>	x"03000001",
		2445 =>	x"00010000",
		2446 =>	x"03000000",
		2447 =>	x"00000303",
		2448 =>	x"03000001",
		2449 =>	x"00010000",
		2450 =>	x"03030300",
		2451 =>	x"00000303",
		2452 =>	x"03000203",
		2453 =>	x"02030200",
		2454 =>	x"03030300",
		2455 =>	x"00000303",
		2456 =>	x"03000202",
		2457 =>	x"02020200",
		2458 =>	x"03030300",
		2459 =>	x"00000003",
		2460 =>	x"03030302",
		2461 =>	x"02020303",
		2462 =>	x"03030000",
		2463 =>	x"00000000",
		2464 =>	x"03030301",
		2465 =>	x"01010303",
		2466 =>	x"03000000",
		2467 =>	x"00000003",
		2468 =>	x"03030301",
		2469 =>	x"01010303",
		2470 =>	x"03030000",
		2471 =>	x"00000303",
		2472 =>	x"03030302",
		2473 =>	x"02020303",
		2474 =>	x"03030300",
		2475 =>	x"00000003",
		2476 =>	x"03030001",
		2477 =>	x"01010003",
		2478 =>	x"03030000",
		2479 =>	x"00000000",
		2480 =>	x"00030000",
		2481 =>	x"00000003",
		2482 =>	x"00000000",
		2483 =>	x"00000000",
		2484 =>	x"00000000",
		2485 =>	x"00000000",
		2486 =>	x"00000000",
		2487 =>	x"00000000",
		2488 =>	x"00000000",
		2489 =>	x"00000000",
		2490 =>	x"00000000",
		2491 =>	x"00000000",
		2492 =>	x"00000000",
		2493 =>	x"00000000",
		2494 =>	x"00000000",
		2495 =>	x"00000000", -- IMG_16x16_muva3_12_skupljeno
		2496 =>	x"00000000",
		2497 =>	x"00000000",
		2498 =>	x"00000000",
		2499 =>	x"00000000",
		2500 =>	x"00000000",
		2501 =>	x"00000000",
		2502 =>	x"00000000",
		2503 =>	x"00000000",
		2504 =>	x"00000000",
		2505 =>	x"00000000",
		2506 =>	x"00000000",
		2507 =>	x"00000003",
		2508 =>	x"00000000",
		2509 =>	x"00000003",
		2510 =>	x"00000000",
		2511 =>	x"00000003",
		2512 =>	x"00000100",
		2513 =>	x"01000003",
		2514 =>	x"00000000",
		2515 =>	x"00000003",
		2516 =>	x"00020302",
		2517 =>	x"03020003",
		2518 =>	x"00000000",
		2519 =>	x"00000003",
		2520 =>	x"00020202",
		2521 =>	x"02020003",
		2522 =>	x"00000000",
		2523 =>	x"00000003",
		2524 =>	x"03030202",
		2525 =>	x"02030303",
		2526 =>	x"00000000",
		2527 =>	x"00000000",
		2528 =>	x"00030101",
		2529 =>	x"01030000",
		2530 =>	x"00000000",
		2531 =>	x"00000003",
		2532 =>	x"03030101",
		2533 =>	x"01030303",
		2534 =>	x"00000000",
		2535 =>	x"00000003",
		2536 =>	x"03030202",
		2537 =>	x"02030303",
		2538 =>	x"00000000",
		2539 =>	x"00000003",
		2540 =>	x"03000101",
		2541 =>	x"01000303",
		2542 =>	x"00000000",
		2543 =>	x"00000003",
		2544 =>	x"03000001",
		2545 =>	x"00000303",
		2546 =>	x"00000000",
		2547 =>	x"00000000",
		2548 =>	x"00000000",
		2549 =>	x"00000000",
		2550 =>	x"00000000",
		2551 =>	x"00000000",
		2552 =>	x"00000000",
		2553 =>	x"00000000",
		2554 =>	x"00000000",
		2555 =>	x"00000000",
		2556 =>	x"00000000",
		2557 =>	x"00000000",
		2558 =>	x"00000000",
		2559 =>	x"00000000", -- IMG_16x16_muva3_9
		2560 =>	x"00000000",
		2561 =>	x"00000000",
		2562 =>	x"00000000",
		2563 =>	x"00000000",
		2564 =>	x"00000000",
		2565 =>	x"00000000",
		2566 =>	x"00000000",
		2567 =>	x"00000000",
		2568 =>	x"03030300",
		2569 =>	x"00000300",
		2570 =>	x"00000000",
		2571 =>	x"00000000",
		2572 =>	x"03030303",
		2573 =>	x"00030303",
		2574 =>	x"00000000",
		2575 =>	x"00000003",
		2576 =>	x"03030303",
		2577 =>	x"03030303",
		2578 =>	x"00000000",
		2579 =>	x"00000000",
		2580 =>	x"00000003",
		2581 =>	x"03030303",
		2582 =>	x"03000000",
		2583 =>	x"00000000",
		2584 =>	x"00020203",
		2585 =>	x"03030300",
		2586 =>	x"00000000",
		2587 =>	x"00000001",
		2588 =>	x"01030202",
		2589 =>	x"01010201",
		2590 =>	x"00000000",
		2591 =>	x"00000000",
		2592 =>	x"00020202",
		2593 =>	x"01010201",
		2594 =>	x"00000000",
		2595 =>	x"00000001",
		2596 =>	x"01030202",
		2597 =>	x"01010201",
		2598 =>	x"00000000",
		2599 =>	x"00000000",
		2600 =>	x"00020203",
		2601 =>	x"03030300",
		2602 =>	x"00000000",
		2603 =>	x"00000000",
		2604 =>	x"00000003",
		2605 =>	x"03030303",
		2606 =>	x"03000000",
		2607 =>	x"00000003",
		2608 =>	x"03030303",
		2609 =>	x"03030303",
		2610 =>	x"00000000",
		2611 =>	x"00000000",
		2612 =>	x"03030303",
		2613 =>	x"00030303",
		2614 =>	x"00000000",
		2615 =>	x"00000000",
		2616 =>	x"03030300",
		2617 =>	x"00000300",
		2618 =>	x"00000000",
		2619 =>	x"00000000",
		2620 =>	x"00000000",
		2621 =>	x"00000000",
		2622 =>	x"00000000",
		2623 =>	x"00000000", -- IMG_16x16_muva3_poal10
		2624 =>	x"00000000",
		2625 =>	x"00000000",
		2626 =>	x"00000000",
		2627 =>	x"00000000",
		2628 =>	x"00000000",
		2629 =>	x"00000000",
		2630 =>	x"00000000",
		2631 =>	x"00000000",
		2632 =>	x"03030300",
		2633 =>	x"00000000",
		2634 =>	x"00000000",
		2635 =>	x"00000000",
		2636 =>	x"00000003",
		2637 =>	x"03000000",
		2638 =>	x"00000000",
		2639 =>	x"00000000",
		2640 =>	x"00000200",
		2641 =>	x"03000303",
		2642 =>	x"03030000",
		2643 =>	x"00000000",
		2644 =>	x"00010301",
		2645 =>	x"03030303",
		2646 =>	x"03030000",
		2647 =>	x"00000000",
		2648 =>	x"00020101",
		2649 =>	x"02020303",
		2650 =>	x"00000000",
		2651 =>	x"00000000",
		2652 =>	x"01030101",
		2653 =>	x"02020101",
		2654 =>	x"00000000",
		2655 =>	x"00000000",
		2656 =>	x"00020101",
		2657 =>	x"02020101",
		2658 =>	x"01000000",
		2659 =>	x"00000000",
		2660 =>	x"00000103",
		2661 =>	x"03020101",
		2662 =>	x"00000000",
		2663 =>	x"00000303",
		2664 =>	x"03000300",
		2665 =>	x"03030300",
		2666 =>	x"00000000",
		2667 =>	x"00000000",
		2668 =>	x"00030300",
		2669 =>	x"03030303",
		2670 =>	x"00000000",
		2671 =>	x"00000000",
		2672 =>	x"00000000",
		2673 =>	x"00000303",
		2674 =>	x"00000000",
		2675 =>	x"00000000",
		2676 =>	x"00000000",
		2677 =>	x"00000000",
		2678 =>	x"00000000",
		2679 =>	x"00000000",
		2680 =>	x"00000000",
		2681 =>	x"00000000",
		2682 =>	x"00000000",
		2683 =>	x"00000000",
		2684 =>	x"00000000",
		2685 =>	x"00000000",
		2686 =>	x"00000000",
		2687 =>	x"00000000", -- IMG_16x16_muva3_pola11
		2688 =>	x"00000000",
		2689 =>	x"00000000",
		2690 =>	x"00000000",
		2691 =>	x"00000000",
		2692 =>	x"00000000",
		2693 =>	x"00000000",
		2694 =>	x"00000000",
		2695 =>	x"00000000",
		2696 =>	x"00000003",
		2697 =>	x"03000000",
		2698 =>	x"00000000",
		2699 =>	x"00000000",
		2700 =>	x"00000000",
		2701 =>	x"03030000",
		2702 =>	x"00000000",
		2703 =>	x"00000000",
		2704 =>	x"00010002",
		2705 =>	x"00030300",
		2706 =>	x"00000000",
		2707 =>	x"00000000",
		2708 =>	x"01000302",
		2709 =>	x"00030000",
		2710 =>	x"00000000",
		2711 =>	x"00000000",
		2712 =>	x"00030202",
		2713 =>	x"02030003",
		2714 =>	x"03000000",
		2715 =>	x"00000300",
		2716 =>	x"02020202",
		2717 =>	x"01010303",
		2718 =>	x"03030000",
		2719 =>	x"00000303",
		2720 =>	x"00000201",
		2721 =>	x"01010200",
		2722 =>	x"03030000",
		2723 =>	x"00000003",
		2724 =>	x"03030301",
		2725 =>	x"01020201",
		2726 =>	x"00000000",
		2727 =>	x"00000000",
		2728 =>	x"03000003",
		2729 =>	x"02020101",
		2730 =>	x"00000000",
		2731 =>	x"00000000",
		2732 =>	x"00000303",
		2733 =>	x"00010101",
		2734 =>	x"00000000",
		2735 =>	x"00000000",
		2736 =>	x"00000303",
		2737 =>	x"03000000",
		2738 =>	x"00000000",
		2739 =>	x"00000000",
		2740 =>	x"00000003",
		2741 =>	x"03000000",
		2742 =>	x"00000000",
		2743 =>	x"00000000",
		2744 =>	x"00000000",
		2745 =>	x"00000000",
		2746 =>	x"00000000",
		2747 =>	x"00000000",
		2748 =>	x"00000000",
		2749 =>	x"00000000",
		2750 =>	x"00000000",
		2751 =>	x"00000000", -- IMG_16x16_muva3_pola12
		2752 =>	x"00000000",
		2753 =>	x"00000000",
		2754 =>	x"00000000",
		2755 =>	x"00000000",
		2756 =>	x"00000000",
		2757 =>	x"00000000",
		2758 =>	x"00000000",
		2759 =>	x"00000000",
		2760 =>	x"00000000",
		2761 =>	x"00000003",
		2762 =>	x"00000000",
		2763 =>	x"00000000",
		2764 =>	x"00000000",
		2765 =>	x"00000003",
		2766 =>	x"00000000",
		2767 =>	x"00000003",
		2768 =>	x"00000000",
		2769 =>	x"01000003",
		2770 =>	x"00000000",
		2771 =>	x"00000003",
		2772 =>	x"00000102",
		2773 =>	x"03020000",
		2774 =>	x"03000000",
		2775 =>	x"00000003",
		2776 =>	x"00020301",
		2777 =>	x"01010103",
		2778 =>	x"03000000",
		2779 =>	x"00000000",
		2780 =>	x"03000101",
		2781 =>	x"01010300",
		2782 =>	x"00000000",
		2783 =>	x"00000000",
		2784 =>	x"03030302",
		2785 =>	x"02020303",
		2786 =>	x"03000000",
		2787 =>	x"00000000",
		2788 =>	x"00000302",
		2789 =>	x"02020203",
		2790 =>	x"03000000",
		2791 =>	x"00000000",
		2792 =>	x"00030303",
		2793 =>	x"01010103",
		2794 =>	x"03030000",
		2795 =>	x"00000000",
		2796 =>	x"00030303",
		2797 =>	x"01010100",
		2798 =>	x"03030000",
		2799 =>	x"00000000",
		2800 =>	x"00030300",
		2801 =>	x"00010000",
		2802 =>	x"00000000",
		2803 =>	x"00000000",
		2804 =>	x"00030300",
		2805 =>	x"00000000",
		2806 =>	x"00000000",
		2807 =>	x"00000000",
		2808 =>	x"00000000",
		2809 =>	x"00000000",
		2810 =>	x"00000000",
		2811 =>	x"00000000",
		2812 =>	x"00000000",
		2813 =>	x"00000000",
		2814 =>	x"00000000",
		2815 =>	x"00000000", -- IMG_16x16_muva4_10
		2816 =>	x"00000000",
		2817 =>	x"00000000",
		2818 =>	x"00000000",
		2819 =>	x"00000000",
		2820 =>	x"00000100",
		2821 =>	x"00000000",
		2822 =>	x"00000000",
		2823 =>	x"00000000",
		2824 =>	x"00000100",
		2825 =>	x"00000000",
		2826 =>	x"00000000",
		2827 =>	x"00000000",
		2828 =>	x"00000001",
		2829 =>	x"00000000",
		2830 =>	x"01010000",
		2831 =>	x"00000000",
		2832 =>	x"000B0300",
		2833 =>	x"01010101",
		2834 =>	x"01010100",
		2835 =>	x"0000000B",
		2836 =>	x"0B03030B",
		2837 =>	x"01010101",
		2838 =>	x"01010100",
		2839 =>	x"00000000",
		2840 =>	x"030B0B0B",
		2841 =>	x"03010001",
		2842 =>	x"00010000",
		2843 =>	x"0000000B",
		2844 =>	x"030B0B0B",
		2845 =>	x"03030B00",
		2846 =>	x"00000000",
		2847 =>	x"00000000",
		2848 =>	x"010B0B03",
		2849 =>	x"030B0B03",
		2850 =>	x"00000000",
		2851 =>	x"00000101",
		2852 =>	x"00010101",
		2853 =>	x"030B0303",
		2854 =>	x"00000000",
		2855 =>	x"00000000",
		2856 =>	x"00000101",
		2857 =>	x"00000300",
		2858 =>	x"00000000",
		2859 =>	x"00000000",
		2860 =>	x"00000101",
		2861 =>	x"01000000",
		2862 =>	x"00000000",
		2863 =>	x"00000000",
		2864 =>	x"00000101",
		2865 =>	x"01000000",
		2866 =>	x"00000000",
		2867 =>	x"00000000",
		2868 =>	x"00000101",
		2869 =>	x"01010000",
		2870 =>	x"00000000",
		2871 =>	x"00000000",
		2872 =>	x"00000001",
		2873 =>	x"01010000",
		2874 =>	x"00000000",
		2875 =>	x"00000000",
		2876 =>	x"00000000",
		2877 =>	x"00000000",
		2878 =>	x"00000000",
		2879 =>	x"00000000", -- IMG_16x16_muva4_11
		2880 =>	x"00000000",
		2881 =>	x"00000000",
		2882 =>	x"00000000",
		2883 =>	x"00000000",
		2884 =>	x"00000000",
		2885 =>	x"00010000",
		2886 =>	x"00000000",
		2887 =>	x"00000000",
		2888 =>	x"000B000B",
		2889 =>	x"00010000",
		2890 =>	x"00000000",
		2891 =>	x"00000000",
		2892 =>	x"000B0303",
		2893 =>	x"01000000",
		2894 =>	x"00000000",
		2895 =>	x"00000000",
		2896 =>	x"0B030B0B",
		2897 =>	x"0B010000",
		2898 =>	x"00000000",
		2899 =>	x"00010100",
		2900 =>	x"03030B0B",
		2901 =>	x"0B010101",
		2902 =>	x"01010000",
		2903 =>	x"00000001",
		2904 =>	x"000B0B0B",
		2905 =>	x"03010101",
		2906 =>	x"01010100",
		2907 =>	x"00000000",
		2908 =>	x"01010303",
		2909 =>	x"03030001",
		2910 =>	x"01010100",
		2911 =>	x"00000000",
		2912 =>	x"01010103",
		2913 =>	x"0B0B0000",
		2914 =>	x"00010100",
		2915 =>	x"00000000",
		2916 =>	x"0101000B",
		2917 =>	x"0B030300",
		2918 =>	x"00000000",
		2919 =>	x"00000000",
		2920 =>	x"01010100",
		2921 =>	x"03030000",
		2922 =>	x"00000000",
		2923 =>	x"00000001",
		2924 =>	x"01010000",
		2925 =>	x"00000000",
		2926 =>	x"00000000",
		2927 =>	x"00000001",
		2928 =>	x"01010100",
		2929 =>	x"00000000",
		2930 =>	x"00000000",
		2931 =>	x"00000000",
		2932 =>	x"01010000",
		2933 =>	x"00000000",
		2934 =>	x"00000000",
		2935 =>	x"00000000",
		2936 =>	x"00000000",
		2937 =>	x"00000000",
		2938 =>	x"00000000",
		2939 =>	x"00000000",
		2940 =>	x"00000000",
		2941 =>	x"00000000",
		2942 =>	x"00000000",
		2943 =>	x"00000000", -- IMG_16x16_muva4_12_rasireno
		2944 =>	x"00000000",
		2945 =>	x"00000000",
		2946 =>	x"00000000",
		2947 =>	x"00000000",
		2948 =>	x"00000000",
		2949 =>	x"00000000",
		2950 =>	x"00000000",
		2951 =>	x"00000000",
		2952 =>	x"00000000",
		2953 =>	x"00000000",
		2954 =>	x"00000000",
		2955 =>	x"00000001",
		2956 =>	x"00000000",
		2957 =>	x"0B000000",
		2958 =>	x"00010000",
		2959 =>	x"00000000",
		2960 =>	x"01000B03",
		2961 =>	x"0B030B00",
		2962 =>	x"01000000",
		2963 =>	x"00000000",
		2964 =>	x"00010303",
		2965 =>	x"0B030301",
		2966 =>	x"00000000",
		2967 =>	x"00000000",
		2968 =>	x"00000B0B",
		2969 =>	x"0B0B0B00",
		2970 =>	x"00000000",
		2971 =>	x"00000000",
		2972 =>	x"0001010B",
		2973 =>	x"0B0B0101",
		2974 =>	x"00000000",
		2975 =>	x"00000000",
		2976 =>	x"01010103",
		2977 =>	x"03030101",
		2978 =>	x"01000000",
		2979 =>	x"00000001",
		2980 =>	x"01010003",
		2981 =>	x"03030001",
		2982 =>	x"01010000",
		2983 =>	x"00000101",
		2984 =>	x"0101000B",
		2985 =>	x"0B0B0001",
		2986 =>	x"01010100",
		2987 =>	x"00000101",
		2988 =>	x"01000003",
		2989 =>	x"03030000",
		2990 =>	x"01010100",
		2991 =>	x"00000101",
		2992 =>	x"01000000",
		2993 =>	x"03000000",
		2994 =>	x"01010100",
		2995 =>	x"00000000",
		2996 =>	x"00000000",
		2997 =>	x"00000000",
		2998 =>	x"00000000",
		2999 =>	x"00000000",
		3000 =>	x"00000000",
		3001 =>	x"00000000",
		3002 =>	x"00000000",
		3003 =>	x"00000000",
		3004 =>	x"00000000",
		3005 =>	x"00000000",
		3006 =>	x"00000000",
		3007 =>	x"00000000", -- IMG_16x16_muva4_12_skupljeno
		3008 =>	x"00000000",
		3009 =>	x"00000000",
		3010 =>	x"00000000",
		3011 =>	x"00000000",
		3012 =>	x"00000000",
		3013 =>	x"00000000",
		3014 =>	x"00000000",
		3015 =>	x"00000000",
		3016 =>	x"00000000",
		3017 =>	x"00000000",
		3018 =>	x"00000000",
		3019 =>	x"00000000",
		3020 =>	x"01000000",
		3021 =>	x"0B000000",
		3022 =>	x"01000000",
		3023 =>	x"00000000",
		3024 =>	x"01000B03",
		3025 =>	x"0B030B00",
		3026 =>	x"01000000",
		3027 =>	x"00000000",
		3028 =>	x"00010303",
		3029 =>	x"0B030301",
		3030 =>	x"00000000",
		3031 =>	x"00000000",
		3032 =>	x"00000B0B",
		3033 =>	x"0B0B0B00",
		3034 =>	x"00000000",
		3035 =>	x"00000000",
		3036 =>	x"0001010B",
		3037 =>	x"0B0B0101",
		3038 =>	x"00000000",
		3039 =>	x"00000000",
		3040 =>	x"00010103",
		3041 =>	x"03030101",
		3042 =>	x"00000000",
		3043 =>	x"00000000",
		3044 =>	x"01010003",
		3045 =>	x"03030001",
		3046 =>	x"01000000",
		3047 =>	x"00000000",
		3048 =>	x"0101000B",
		3049 =>	x"0B0B0001",
		3050 =>	x"01000000",
		3051 =>	x"00000000",
		3052 =>	x"01010003",
		3053 =>	x"03030001",
		3054 =>	x"01000000",
		3055 =>	x"00000000",
		3056 =>	x"01010000",
		3057 =>	x"03000001",
		3058 =>	x"01000000",
		3059 =>	x"00000000",
		3060 =>	x"00000000",
		3061 =>	x"00000000",
		3062 =>	x"00000000",
		3063 =>	x"00000000",
		3064 =>	x"00000000",
		3065 =>	x"00000000",
		3066 =>	x"00000000",
		3067 =>	x"00000000",
		3068 =>	x"00000000",
		3069 =>	x"00000000",
		3070 =>	x"00000000",
		3071 =>	x"00000000", -- IMG_16x16_muva4_9
		3072 =>	x"00000000",
		3073 =>	x"00000000",
		3074 =>	x"00000000",
		3075 =>	x"00000000",
		3076 =>	x"00000000",
		3077 =>	x"00000000",
		3078 =>	x"00000000",
		3079 =>	x"00000000",
		3080 =>	x"00000000",
		3081 =>	x"00000101",
		3082 =>	x"01000000",
		3083 =>	x"00000001",
		3084 =>	x"00000000",
		3085 =>	x"00010101",
		3086 =>	x"01000000",
		3087 =>	x"00000000",
		3088 =>	x"01000000",
		3089 =>	x"01010101",
		3090 =>	x"01000000",
		3091 =>	x"00000000",
		3092 =>	x"00010001",
		3093 =>	x"01010100",
		3094 =>	x"00000000",
		3095 =>	x"00000000",
		3096 =>	x"0B030B01",
		3097 =>	x"01000000",
		3098 =>	x"00000000",
		3099 =>	x"00000000",
		3100 =>	x"03030B0B",
		3101 =>	x"03030B03",
		3102 =>	x"00000000",
		3103 =>	x"0000000B",
		3104 =>	x"0B0B0B0B",
		3105 =>	x"03030B03",
		3106 =>	x"03000000",
		3107 =>	x"00000000",
		3108 =>	x"03030B0B",
		3109 =>	x"03030B03",
		3110 =>	x"00000000",
		3111 =>	x"00000000",
		3112 =>	x"0B030B01",
		3113 =>	x"01000000",
		3114 =>	x"00000000",
		3115 =>	x"00000000",
		3116 =>	x"00010001",
		3117 =>	x"01010100",
		3118 =>	x"00000000",
		3119 =>	x"00000000",
		3120 =>	x"01000000",
		3121 =>	x"01010101",
		3122 =>	x"01000000",
		3123 =>	x"00000001",
		3124 =>	x"00000000",
		3125 =>	x"00010101",
		3126 =>	x"01000000",
		3127 =>	x"00000000",
		3128 =>	x"00000000",
		3129 =>	x"00000101",
		3130 =>	x"01000000",
		3131 =>	x"00000000",
		3132 =>	x"00000000",
		3133 =>	x"00000000",
		3134 =>	x"00000000",
		3135 =>	x"00000000", -- IMG_16x16_muva4_pola10
		3136 =>	x"00000000",
		3137 =>	x"00000000",
		3138 =>	x"00000000",
		3139 =>	x"00000000",
		3140 =>	x"00000000",
		3141 =>	x"00000000",
		3142 =>	x"00000000",
		3143 =>	x"00000000",
		3144 =>	x"00000000",
		3145 =>	x"00000000",
		3146 =>	x"00000000",
		3147 =>	x"00000000",
		3148 =>	x"00010000",
		3149 =>	x"00000000",
		3150 =>	x"00000000",
		3151 =>	x"00000000",
		3152 =>	x"00000100",
		3153 =>	x"00000000",
		3154 =>	x"00000000",
		3155 =>	x"00000000",
		3156 =>	x"000B0100",
		3157 =>	x"01010101",
		3158 =>	x"01010000",
		3159 =>	x"00000000",
		3160 =>	x"03030B0B",
		3161 =>	x"01010101",
		3162 =>	x"01010000",
		3163 =>	x"0000000B",
		3164 =>	x"0B0B0B0B",
		3165 =>	x"03030000",
		3166 =>	x"00000000",
		3167 =>	x"00000000",
		3168 =>	x"03030B0B",
		3169 =>	x"03030B03",
		3170 =>	x"00000000",
		3171 =>	x"00000000",
		3172 =>	x"0B030B0B",
		3173 =>	x"03030B03",
		3174 =>	x"03000000",
		3175 =>	x"00000000",
		3176 =>	x"01000101",
		3177 =>	x"00030B03",
		3178 =>	x"00000000",
		3179 =>	x"00000101",
		3180 =>	x"00000101",
		3181 =>	x"01000000",
		3182 =>	x"00000000",
		3183 =>	x"00000000",
		3184 =>	x"00000000",
		3185 =>	x"01010101",
		3186 =>	x"00000000",
		3187 =>	x"00000000",
		3188 =>	x"00000000",
		3189 =>	x"00010101",
		3190 =>	x"00000000",
		3191 =>	x"00000000",
		3192 =>	x"00000000",
		3193 =>	x"00000000",
		3194 =>	x"00000000",
		3195 =>	x"00000000",
		3196 =>	x"00000000",
		3197 =>	x"00000000",
		3198 =>	x"00000000",
		3199 =>	x"00000000", -- IMG_16x16_muva4_pola11
		3200 =>	x"00000000",
		3201 =>	x"00000000",
		3202 =>	x"00000000",
		3203 =>	x"00000000",
		3204 =>	x"00000000",
		3205 =>	x"00000000",
		3206 =>	x"00000000",
		3207 =>	x"00000000",
		3208 =>	x"00000001",
		3209 =>	x"00000000",
		3210 =>	x"00000000",
		3211 =>	x"00000000",
		3212 =>	x"00000000",
		3213 =>	x"01000000",
		3214 =>	x"00000000",
		3215 =>	x"00000000",
		3216 =>	x"0B00030B",
		3217 =>	x"01000000",
		3218 =>	x"00000000",
		3219 =>	x"00000000",
		3220 =>	x"000B0303",
		3221 =>	x"0B010000",
		3222 =>	x"00000000",
		3223 =>	x"00000000",
		3224 =>	x"03030B0B",
		3225 =>	x"0B010101",
		3226 =>	x"01000000",
		3227 =>	x"00000100",
		3228 =>	x"0B030B0B",
		3229 =>	x"0B030B01",
		3230 =>	x"01010000",
		3231 =>	x"00000001",
		3232 =>	x"010B0B0B",
		3233 =>	x"03030B01",
		3234 =>	x"01010100",
		3235 =>	x"00000000",
		3236 =>	x"00010103",
		3237 =>	x"030B0B03",
		3238 =>	x"00010000",
		3239 =>	x"00000000",
		3240 =>	x"0000010B",
		3241 =>	x"0B0B0300",
		3242 =>	x"00000000",
		3243 =>	x"00000000",
		3244 =>	x"00000101",
		3245 =>	x"01030003",
		3246 =>	x"00000000",
		3247 =>	x"00000000",
		3248 =>	x"00000101",
		3249 =>	x"01000000",
		3250 =>	x"00000000",
		3251 =>	x"00000000",
		3252 =>	x"00000001",
		3253 =>	x"01010000",
		3254 =>	x"00000000",
		3255 =>	x"00000000",
		3256 =>	x"00000000",
		3257 =>	x"01000000",
		3258 =>	x"00000000",
		3259 =>	x"00000000",
		3260 =>	x"00000000",
		3261 =>	x"00000000",
		3262 =>	x"00000000",
		3263 =>	x"00000000", -- IMG_16x16_muva4_pola12
		3264 =>	x"00000000",
		3265 =>	x"00000000",
		3266 =>	x"00000000",
		3267 =>	x"00000000",
		3268 =>	x"00000000",
		3269 =>	x"00000000",
		3270 =>	x"00000000",
		3271 =>	x"00000000",
		3272 =>	x"00000000",
		3273 =>	x"00000100",
		3274 =>	x"00000000",
		3275 =>	x"00000000",
		3276 =>	x"00000B00",
		3277 =>	x"00000100",
		3278 =>	x"00000000",
		3279 =>	x"00000000",
		3280 =>	x"00030B03",
		3281 =>	x"0B010000",
		3282 =>	x"00000000",
		3283 =>	x"00000100",
		3284 =>	x"0B030B03",
		3285 =>	x"03000000",
		3286 =>	x"00000000",
		3287 =>	x"00000001",
		3288 =>	x"010B0B0B",
		3289 =>	x"0B010100",
		3290 =>	x"00000000",
		3291 =>	x"00000000",
		3292 =>	x"000B0B0B",
		3293 =>	x"0B010100",
		3294 =>	x"00000000",
		3295 =>	x"00000000",
		3296 =>	x"01010303",
		3297 =>	x"03000101",
		3298 =>	x"00000000",
		3299 =>	x"00000000",
		3300 =>	x"01010303",
		3301 =>	x"03030001",
		3302 =>	x"01000000",
		3303 =>	x"00000000",
		3304 =>	x"0101000B",
		3305 =>	x"0B0B0001",
		3306 =>	x"01000000",
		3307 =>	x"00000000",
		3308 =>	x"01010003",
		3309 =>	x"03030001",
		3310 =>	x"01000000",
		3311 =>	x"00000000",
		3312 =>	x"01010000",
		3313 =>	x"03000000",
		3314 =>	x"00000000",
		3315 =>	x"00000000",
		3316 =>	x"01010000",
		3317 =>	x"00000000",
		3318 =>	x"00000000",
		3319 =>	x"00000000",
		3320 =>	x"00000000",
		3321 =>	x"00000000",
		3322 =>	x"00000000",
		3323 =>	x"00000000",
		3324 =>	x"00000000",
		3325 =>	x"00000000",
		3326 =>	x"00000000",
		3327 =>	x"00000000", -- IMG_16x16_muva5_10
		3328 =>	x"00000000",
		3329 =>	x"00000000",
		3330 =>	x"00000000",
		3331 =>	x"00000000",
		3332 =>	x"00000000",
		3333 =>	x"00010000",
		3334 =>	x"00000000",
		3335 =>	x"00000000",
		3336 =>	x"00000000",
		3337 =>	x"00010000",
		3338 =>	x"00000000",
		3339 =>	x"00000000",
		3340 =>	x"00000000",
		3341 =>	x"01010202",
		3342 =>	x"00000000",
		3343 =>	x"00000000",
		3344 =>	x"03000000",
		3345 =>	x"01010200",
		3346 =>	x"00000000",
		3347 =>	x"00000000",
		3348 =>	x"03030001",
		3349 =>	x"01020202",
		3350 =>	x"00000000",
		3351 =>	x"00000000",
		3352 =>	x"01000001",
		3353 =>	x"01020200",
		3354 =>	x"00000000",
		3355 =>	x"00000303",
		3356 =>	x"03010101",
		3357 =>	x"02020000",
		3358 =>	x"00000000",
		3359 =>	x"00000000",
		3360 =>	x"00000101",
		3361 =>	x"01000000",
		3362 =>	x"00000000",
		3363 =>	x"00000000",
		3364 =>	x"00010102",
		3365 =>	x"00010100",
		3366 =>	x"00000000",
		3367 =>	x"00000000",
		3368 =>	x"01010202",
		3369 =>	x"00000101",
		3370 =>	x"00000000",
		3371 =>	x"00000001",
		3372 =>	x"01010202",
		3373 =>	x"00000000",
		3374 =>	x"01000000",
		3375 =>	x"00000001",
		3376 =>	x"01020200",
		3377 =>	x"00000000",
		3378 =>	x"00010000",
		3379 =>	x"00000101",
		3380 =>	x"02020000",
		3381 =>	x"00000000",
		3382 =>	x"00000000",
		3383 =>	x"00000000",
		3384 =>	x"00000000",
		3385 =>	x"00000000",
		3386 =>	x"00000000",
		3387 =>	x"00000000",
		3388 =>	x"00000000",
		3389 =>	x"00000000",
		3390 =>	x"00000000",
		3391 =>	x"00000000", -- IMG_16x16_muva5_11
		3392 =>	x"00000000",
		3393 =>	x"00000000",
		3394 =>	x"00000000",
		3395 =>	x"00000000",
		3396 =>	x"00000000",
		3397 =>	x"00000000",
		3398 =>	x"00000000",
		3399 =>	x"00000000",
		3400 =>	x"00000003",
		3401 =>	x"00000000",
		3402 =>	x"00010000",
		3403 =>	x"00000000",
		3404 =>	x"00000003",
		3405 =>	x"00000001",
		3406 =>	x"01010000",
		3407 =>	x"00000000",
		3408 =>	x"03030103",
		3409 =>	x"00000101",
		3410 =>	x"01020000",
		3411 =>	x"00000000",
		3412 =>	x"00030001",
		3413 =>	x"00010101",
		3414 =>	x"02020000",
		3415 =>	x"00000000",
		3416 =>	x"00000001",
		3417 =>	x"01010202",
		3418 =>	x"02000000",
		3419 =>	x"00000000",
		3420 =>	x"00010101",
		3421 =>	x"01020202",
		3422 =>	x"00000000",
		3423 =>	x"00000001",
		3424 =>	x"01010102",
		3425 =>	x"01000000",
		3426 =>	x"00000000",
		3427 =>	x"00010101",
		3428 =>	x"01020202",
		3429 =>	x"00010000",
		3430 =>	x"00000000",
		3431 =>	x"00000002",
		3432 =>	x"02020200",
		3433 =>	x"00010100",
		3434 =>	x"00000000",
		3435 =>	x"00000002",
		3436 =>	x"00020000",
		3437 =>	x"00000100",
		3438 =>	x"00000000",
		3439 =>	x"00000000",
		3440 =>	x"00000000",
		3441 =>	x"00000001",
		3442 =>	x"00000000",
		3443 =>	x"00000000",
		3444 =>	x"00000000",
		3445 =>	x"00000000",
		3446 =>	x"01000000",
		3447 =>	x"00000000",
		3448 =>	x"00000000",
		3449 =>	x"00000000",
		3450 =>	x"00000000",
		3451 =>	x"00000000",
		3452 =>	x"00000000",
		3453 =>	x"00000000",
		3454 =>	x"00000000",
		3455 =>	x"00000000", -- IMG_16x16_muva5_12
		3456 =>	x"00000000",
		3457 =>	x"00000000",
		3458 =>	x"00000000",
		3459 =>	x"00000000",
		3460 =>	x"00000000",
		3461 =>	x"00000000",
		3462 =>	x"00000000",
		3463 =>	x"00000000",
		3464 =>	x"00000000",
		3465 =>	x"00000000",
		3466 =>	x"00000000",
		3467 =>	x"00000000",
		3468 =>	x"00000303",
		3469 =>	x"00030300",
		3470 =>	x"00000000",
		3471 =>	x"00000000",
		3472 =>	x"00000003",
		3473 =>	x"01030000",
		3474 =>	x"00000000",
		3475 =>	x"00000000",
		3476 =>	x"00000000",
		3477 =>	x"01000000",
		3478 =>	x"00000000",
		3479 =>	x"00010101",
		3480 =>	x"01010100",
		3481 =>	x"01000101",
		3482 =>	x"01010101",
		3483 =>	x"00000101",
		3484 =>	x"01010101",
		3485 =>	x"01010101",
		3486 =>	x"01010100",
		3487 =>	x"00000202",
		3488 =>	x"02020202",
		3489 =>	x"01020202",
		3490 =>	x"02020200",
		3491 =>	x"00000000",
		3492 =>	x"02020200",
		3493 =>	x"01000202",
		3494 =>	x"02000000",
		3495 =>	x"00000000",
		3496 =>	x"00000000",
		3497 =>	x"01000000",
		3498 =>	x"00000000",
		3499 =>	x"00000000",
		3500 =>	x"00000000",
		3501 =>	x"01000000",
		3502 =>	x"00000000",
		3503 =>	x"00000000",
		3504 =>	x"00000000",
		3505 =>	x"01000000",
		3506 =>	x"00000000",
		3507 =>	x"00000000",
		3508 =>	x"00000000",
		3509 =>	x"01000000",
		3510 =>	x"00000000",
		3511 =>	x"00000000",
		3512 =>	x"00000000",
		3513 =>	x"01000000",
		3514 =>	x"00000000",
		3515 =>	x"00000000",
		3516 =>	x"00000000",
		3517 =>	x"00000000",
		3518 =>	x"00000000",
		3519 =>	x"00000000", -- IMG_16x16_muva5_9
		3520 =>	x"00000000",
		3521 =>	x"00000000",
		3522 =>	x"00000000",
		3523 =>	x"00000000",
		3524 =>	x"00010000",
		3525 =>	x"00000000",
		3526 =>	x"00000000",
		3527 =>	x"00000000",
		3528 =>	x"00010102",
		3529 =>	x"00000000",
		3530 =>	x"00000000",
		3531 =>	x"00000000",
		3532 =>	x"00010102",
		3533 =>	x"00000000",
		3534 =>	x"00000000",
		3535 =>	x"00000000",
		3536 =>	x"00010102",
		3537 =>	x"02000000",
		3538 =>	x"00000000",
		3539 =>	x"00000000",
		3540 =>	x"00010102",
		3541 =>	x"02000000",
		3542 =>	x"00000000",
		3543 =>	x"00000300",
		3544 =>	x"00010102",
		3545 =>	x"02000000",
		3546 =>	x"00000000",
		3547 =>	x"00000303",
		3548 =>	x"00000102",
		3549 =>	x"00000000",
		3550 =>	x"00000000",
		3551 =>	x"00000001",
		3552 =>	x"01010101",
		3553 =>	x"01010101",
		3554 =>	x"01010000",
		3555 =>	x"00000303",
		3556 =>	x"00000102",
		3557 =>	x"00000000",
		3558 =>	x"00000000",
		3559 =>	x"00000300",
		3560 =>	x"00010102",
		3561 =>	x"02000000",
		3562 =>	x"00000000",
		3563 =>	x"00000000",
		3564 =>	x"00010102",
		3565 =>	x"02000000",
		3566 =>	x"00000000",
		3567 =>	x"00000000",
		3568 =>	x"00010102",
		3569 =>	x"02000000",
		3570 =>	x"00000000",
		3571 =>	x"00000000",
		3572 =>	x"00010102",
		3573 =>	x"00000000",
		3574 =>	x"00000000",
		3575 =>	x"00000000",
		3576 =>	x"00010102",
		3577 =>	x"00000000",
		3578 =>	x"00000000",
		3579 =>	x"00000000",
		3580 =>	x"00010000",
		3581 =>	x"00000000",
		3582 =>	x"00000000",
		3583 =>	x"00000000", -- IMG_16x16_muva5_pola10
		3584 =>	x"00000000",
		3585 =>	x"00000000",
		3586 =>	x"00000000",
		3587 =>	x"00000000",
		3588 =>	x"00000001",
		3589 =>	x"00000000",
		3590 =>	x"00000000",
		3591 =>	x"00000000",
		3592 =>	x"00000001",
		3593 =>	x"01000000",
		3594 =>	x"00000000",
		3595 =>	x"00000000",
		3596 =>	x"00000001",
		3597 =>	x"01020000",
		3598 =>	x"00000000",
		3599 =>	x"00000000",
		3600 =>	x"00000101",
		3601 =>	x"01020000",
		3602 =>	x"00000000",
		3603 =>	x"00000003",
		3604 =>	x"00000101",
		3605 =>	x"02020000",
		3606 =>	x"00000000",
		3607 =>	x"00000003",
		3608 =>	x"03000101",
		3609 =>	x"02020000",
		3610 =>	x"00000000",
		3611 =>	x"00000000",
		3612 =>	x"01000001",
		3613 =>	x"02020000",
		3614 =>	x"00000000",
		3615 =>	x"00000303",
		3616 =>	x"00010101",
		3617 =>	x"01000000",
		3618 =>	x"00000000",
		3619 =>	x"00000300",
		3620 =>	x"00000102",
		3621 =>	x"00010101",
		3622 =>	x"00000000",
		3623 =>	x"00000000",
		3624 =>	x"00010102",
		3625 =>	x"00000000",
		3626 =>	x"01010000",
		3627 =>	x"00000000",
		3628 =>	x"00010202",
		3629 =>	x"02000000",
		3630 =>	x"00000000",
		3631 =>	x"00000000",
		3632 =>	x"01010202",
		3633 =>	x"00000000",
		3634 =>	x"00000000",
		3635 =>	x"00000000",
		3636 =>	x"01010200",
		3637 =>	x"00000000",
		3638 =>	x"00000000",
		3639 =>	x"00000001",
		3640 =>	x"01020200",
		3641 =>	x"00000000",
		3642 =>	x"00000000",
		3643 =>	x"00000000",
		3644 =>	x"00000000",
		3645 =>	x"00000000",
		3646 =>	x"00000000",
		3647 =>	x"00000000", -- IMG_16x16_muva5_pola11
		3648 =>	x"00000000",
		3649 =>	x"00000000",
		3650 =>	x"00000000",
		3651 =>	x"00000000",
		3652 =>	x"00000000",
		3653 =>	x"00000001",
		3654 =>	x"00000000",
		3655 =>	x"00000000",
		3656 =>	x"00000000",
		3657 =>	x"00000101",
		3658 =>	x"00000000",
		3659 =>	x"00000000",
		3660 =>	x"00030000",
		3661 =>	x"00010101",
		3662 =>	x"02000000",
		3663 =>	x"00000000",
		3664 =>	x"00030300",
		3665 =>	x"00010102",
		3666 =>	x"02000000",
		3667 =>	x"00000003",
		3668 =>	x"03010000",
		3669 =>	x"01010202",
		3670 =>	x"00000000",
		3671 =>	x"00000000",
		3672 =>	x"03000100",
		3673 =>	x"01020202",
		3674 =>	x"00000000",
		3675 =>	x"00000000",
		3676 =>	x"00000001",
		3677 =>	x"02020200",
		3678 =>	x"00000000",
		3679 =>	x"00000000",
		3680 =>	x"00010102",
		3681 =>	x"01000000",
		3682 =>	x"00000000",
		3683 =>	x"00000001",
		3684 =>	x"01010202",
		3685 =>	x"00010000",
		3686 =>	x"00000000",
		3687 =>	x"00000101",
		3688 =>	x"01020202",
		3689 =>	x"00000100",
		3690 =>	x"00000000",
		3691 =>	x"00010101",
		3692 =>	x"02020200",
		3693 =>	x"00000001",
		3694 =>	x"00000000",
		3695 =>	x"00000002",
		3696 =>	x"02000000",
		3697 =>	x"00000000",
		3698 =>	x"01000000",
		3699 =>	x"00000000",
		3700 =>	x"00000000",
		3701 =>	x"00000000",
		3702 =>	x"00010000",
		3703 =>	x"00000000",
		3704 =>	x"00000000",
		3705 =>	x"00000000",
		3706 =>	x"00000000",
		3707 =>	x"00000000",
		3708 =>	x"00000000",
		3709 =>	x"00000000",
		3710 =>	x"00000000",
		3711 =>	x"00000000", -- IMG_16x16_muva5_pola12
		3712 =>	x"00000000",
		3713 =>	x"00000000",
		3714 =>	x"00000000",
		3715 =>	x"00000000",
		3716 =>	x"00000000",
		3717 =>	x"00000000",
		3718 =>	x"00000000",
		3719 =>	x"00000000",
		3720 =>	x"00000000",
		3721 =>	x"00000000",
		3722 =>	x"00000000",
		3723 =>	x"00000000",
		3724 =>	x"00000003",
		3725 =>	x"03000000",
		3726 =>	x"00000000",
		3727 =>	x"00000000",
		3728 =>	x"03030003",
		3729 =>	x"00000000",
		3730 =>	x"00010000",
		3731 =>	x"00000000",
		3732 =>	x"00030100",
		3733 =>	x"00000001",
		3734 =>	x"01010000",
		3735 =>	x"00000000",
		3736 =>	x"00000001",
		3737 =>	x"00010101",
		3738 =>	x"01020000",
		3739 =>	x"00000001",
		3740 =>	x"01010001",
		3741 =>	x"01010202",
		3742 =>	x"02020000",
		3743 =>	x"01010101",
		3744 =>	x"01010101",
		3745 =>	x"02020202",
		3746 =>	x"00000000",
		3747 =>	x"00010101",
		3748 =>	x"02020201",
		3749 =>	x"00000200",
		3750 =>	x"00000000",
		3751 =>	x"00000202",
		3752 =>	x"02020200",
		3753 =>	x"01000000",
		3754 =>	x"00000000",
		3755 =>	x"00000000",
		3756 =>	x"00000000",
		3757 =>	x"01000000",
		3758 =>	x"00000000",
		3759 =>	x"00000000",
		3760 =>	x"00000000",
		3761 =>	x"01000000",
		3762 =>	x"00000000",
		3763 =>	x"00000000",
		3764 =>	x"00000000",
		3765 =>	x"00010000",
		3766 =>	x"00000000",
		3767 =>	x"00000000",
		3768 =>	x"00000000",
		3769 =>	x"00010000",
		3770 =>	x"00000000",
		3771 =>	x"00000000",
		3772 =>	x"00000000",
		3773 =>	x"00000000",
		3774 =>	x"00000000",
		3775 =>	x"00000000", -- IMG_16x16_muva_10
		3776 =>	x"0C000000",
		3777 =>	x"000C0000",
		3778 =>	x"00000000",
		3779 =>	x"00000000",
		3780 =>	x"0C000000",
		3781 =>	x"0C0C0000",
		3782 =>	x"00000000",
		3783 =>	x"00000C0D",
		3784 =>	x"0D0C000C",
		3785 =>	x"0C0C0C0C",
		3786 =>	x"0C0C0000",
		3787 =>	x"000C0C0C",
		3788 =>	x"0C0C0B0C",
		3789 =>	x"0C0C0D0D",
		3790 =>	x"0D0C0C00",
		3791 =>	x"00000D0D",
		3792 =>	x"0C0B0B0B",
		3793 =>	x"0B0C0C0C",
		3794 =>	x"0D0C0C0C",
		3795 =>	x"00000D0C",
		3796 =>	x"0B0B0B0B",
		3797 =>	x"0D000000",
		3798 =>	x"0C0C0C00",
		3799 =>	x"000C0C00",
		3800 =>	x"0B0B0B0B",
		3801 =>	x"00000000",
		3802 =>	x"00000000",
		3803 =>	x"00000000",
		3804 =>	x"0C0B0B0D",
		3805 =>	x"0D000000",
		3806 =>	x"00000000",
		3807 =>	x"0000000C",
		3808 =>	x"0C0C0C00",
		3809 =>	x"00000000",
		3810 =>	x"00000000",
		3811 =>	x"0000000C",
		3812 =>	x"0C0C0C00",
		3813 =>	x"00000000",
		3814 =>	x"00000000",
		3815 =>	x"0000000C",
		3816 =>	x"0C0C0C0C",
		3817 =>	x"0C000000",
		3818 =>	x"00000000",
		3819 =>	x"00000000",
		3820 =>	x"000C0C0C",
		3821 =>	x"0D0C0C00",
		3822 =>	x"00000000",
		3823 =>	x"00000000",
		3824 =>	x"00000C0D",
		3825 =>	x"0D0C0C00",
		3826 =>	x"00000000",
		3827 =>	x"00000000",
		3828 =>	x"0000000C",
		3829 =>	x"0C0C0C00",
		3830 =>	x"00000000",
		3831 =>	x"00000000",
		3832 =>	x"00000000",
		3833 =>	x"00000000",
		3834 =>	x"00000000",
		3835 =>	x"00000000",
		3836 =>	x"00000000",
		3837 =>	x"00000000",
		3838 =>	x"00000000",
		3839 =>	x"00000000", -- IMG_16x16_muva_11
		3840 =>	x"0C00000C",
		3841 =>	x"00000000",
		3842 =>	x"00000000",
		3843 =>	x"0000000C",
		3844 =>	x"0C0D0D0C",
		3845 =>	x"00000000",
		3846 =>	x"00000000",
		3847 =>	x"0000000D",
		3848 =>	x"0C0D0C00",
		3849 =>	x"000C0C0C",
		3850 =>	x"00000000",
		3851 =>	x"000C0C0D",
		3852 =>	x"0C0C0B0B",
		3853 =>	x"0C0C0C0C",
		3854 =>	x"00000000",
		3855 =>	x"0000000C",
		3856 =>	x"0C0B0B0B",
		3857 =>	x"0B0C0C0C",
		3858 =>	x"0C000000",
		3859 =>	x"00000000",
		3860 =>	x"0B0B0B0B",
		3861 =>	x"0B0C0C0C",
		3862 =>	x"0C0C0000",
		3863 =>	x"0000000C",
		3864 =>	x"0C0B0B0B",
		3865 =>	x"0D00000C",
		3866 =>	x"0C0D0C00",
		3867 =>	x"00000C0C",
		3868 =>	x"0C0B0D00",
		3869 =>	x"0D00000C",
		3870 =>	x"0D0D0C00",
		3871 =>	x"000C0C0C",
		3872 =>	x"0C0C0000",
		3873 =>	x"00000000",
		3874 =>	x"0C0C0C00",
		3875 =>	x"0000000C",
		3876 =>	x"0D0C0000",
		3877 =>	x"00000000",
		3878 =>	x"0C0C0C00",
		3879 =>	x"0000000C",
		3880 =>	x"0D0C0000",
		3881 =>	x"00000000",
		3882 =>	x"00000000",
		3883 =>	x"0000000C",
		3884 =>	x"0D0D0C00",
		3885 =>	x"00000000",
		3886 =>	x"00000000",
		3887 =>	x"0000000C",
		3888 =>	x"0C0C0C00",
		3889 =>	x"00000000",
		3890 =>	x"00000000",
		3891 =>	x"00000000",
		3892 =>	x"0C0C0C00",
		3893 =>	x"00000000",
		3894 =>	x"00000000",
		3895 =>	x"00000000",
		3896 =>	x"000C0000",
		3897 =>	x"00000000",
		3898 =>	x"00000000",
		3899 =>	x"00000000",
		3900 =>	x"00000000",
		3901 =>	x"00000000",
		3902 =>	x"00000000",
		3903 =>	x"00000000", -- IMG_16x16_muva_12_rasireno
		3904 =>	x"0000000C",
		3905 =>	x"000C0000",
		3906 =>	x"00000000",
		3907 =>	x"00000000",
		3908 =>	x"0C0C0D0D",
		3909 =>	x"0C0D0D0C",
		3910 =>	x"0C000000",
		3911 =>	x"00000000",
		3912 =>	x"000C0D0D",
		3913 =>	x"0C0D0D0C",
		3914 =>	x"00000000",
		3915 =>	x"00000000",
		3916 =>	x"00000C0C",
		3917 =>	x"0C0C0C00",
		3918 =>	x"00000000",
		3919 =>	x"00000000",
		3920 =>	x"000C0B0B",
		3921 =>	x"0C0B0B0C",
		3922 =>	x"00000000",
		3923 =>	x"0000000C",
		3924 =>	x"0C0C0B0B",
		3925 =>	x"0B0B0B0C",
		3926 =>	x"0C0C0000",
		3927 =>	x"000C0C0C",
		3928 =>	x"0C0C0B0B",
		3929 =>	x"0B0B0B0C",
		3930 =>	x"0C0C0C0C",
		3931 =>	x"00000C0C",
		3932 =>	x"0C0C0B0B",
		3933 =>	x"0B0B0B0C",
		3934 =>	x"0C0C0C00",
		3935 =>	x"00000C0D",
		3936 =>	x"0C0C000D",
		3937 =>	x"000D000C",
		3938 =>	x"0C0D0C00",
		3939 =>	x"000C0C0D",
		3940 =>	x"0C00000D",
		3941 =>	x"000D0000",
		3942 =>	x"0C0D0C0C",
		3943 =>	x"000C0D0C",
		3944 =>	x"0C000000",
		3945 =>	x"00000000",
		3946 =>	x"0C0C0D0C",
		3947 =>	x"000C0D0D",
		3948 =>	x"0C000000",
		3949 =>	x"00000000",
		3950 =>	x"0C0D0D0C",
		3951 =>	x"000C0D0D",
		3952 =>	x"0C000000",
		3953 =>	x"00000000",
		3954 =>	x"0C0D0D0C",
		3955 =>	x"000C0C0C",
		3956 =>	x"0C000000",
		3957 =>	x"00000000",
		3958 =>	x"0C0C0C0C",
		3959 =>	x"00000C0C",
		3960 =>	x"00000000",
		3961 =>	x"00000000",
		3962 =>	x"000C0C00",
		3963 =>	x"00000000",
		3964 =>	x"00000000",
		3965 =>	x"00000000",
		3966 =>	x"00000000",
		3967 =>	x"00000000", -- IMG_16x16_muva_12_skupljeno
		3968 =>	x"0000000C",
		3969 =>	x"000C0000",
		3970 =>	x"00000000",
		3971 =>	x"00000000",
		3972 =>	x"0C0C0D0D",
		3973 =>	x"0C0D0D0C",
		3974 =>	x"0C000000",
		3975 =>	x"00000000",
		3976 =>	x"000C0D0D",
		3977 =>	x"0C0D0D0C",
		3978 =>	x"00000000",
		3979 =>	x"00000000",
		3980 =>	x"00000C0C",
		3981 =>	x"0C0C0C00",
		3982 =>	x"00000000",
		3983 =>	x"00000000",
		3984 =>	x"0C0C0B0B",
		3985 =>	x"0C0B0B0C",
		3986 =>	x"0C000000",
		3987 =>	x"0000000C",
		3988 =>	x"0C0C0B0B",
		3989 =>	x"0B0B0B0C",
		3990 =>	x"0C0C0000",
		3991 =>	x"000C0C0C",
		3992 =>	x"0C0C0B0B",
		3993 =>	x"0B0B0B0C",
		3994 =>	x"0C0C0C0C",
		3995 =>	x"00000C0C",
		3996 =>	x"0C000B0B",
		3997 =>	x"0B0B0B00",
		3998 =>	x"0C0C0C00",
		3999 =>	x"0000000C",
		4000 =>	x"0C00000D",
		4001 =>	x"000D0000",
		4002 =>	x"0C0C0000",
		4003 =>	x"0000000C",
		4004 =>	x"0C00000D",
		4005 =>	x"000D0000",
		4006 =>	x"0C0C0000",
		4007 =>	x"0000000C",
		4008 =>	x"0C0C0000",
		4009 =>	x"0000000C",
		4010 =>	x"0C0C0000",
		4011 =>	x"00000000",
		4012 =>	x"0C0C0000",
		4013 =>	x"0000000C",
		4014 =>	x"0C000000",
		4015 =>	x"00000000",
		4016 =>	x"000C0C00",
		4017 =>	x"00000C0C",
		4018 =>	x"00000000",
		4019 =>	x"00000000",
		4020 =>	x"00000C0C",
		4021 =>	x"000C0C00",
		4022 =>	x"00000000",
		4023 =>	x"00000000",
		4024 =>	x"0000000C",
		4025 =>	x"000C0000",
		4026 =>	x"00000000",
		4027 =>	x"00000000",
		4028 =>	x"00000000",
		4029 =>	x"00000000",
		4030 =>	x"00000000",
		4031 =>	x"00000000", -- IMG_16x16_muva_9
		4032 =>	x"0000000C",
		4033 =>	x"00000C0C",
		4034 =>	x"0C0C0C00",
		4035 =>	x"00000000",
		4036 =>	x"0000000C",
		4037 =>	x"0C0C0C0D",
		4038 =>	x"0D0D0C0C",
		4039 =>	x"00000000",
		4040 =>	x"00000C0C",
		4041 =>	x"0C0D0D0C",
		4042 =>	x"0D0D0C0C",
		4043 =>	x"00000C00",
		4044 =>	x"00000C0C",
		4045 =>	x"0C0C0C0C",
		4046 =>	x"0C0C0C00",
		4047 =>	x"00000C0C",
		4048 =>	x"000C0C0C",
		4049 =>	x"0C0C0000",
		4050 =>	x"00000000",
		4051 =>	x"00000D0D",
		4052 =>	x"0C0B0B0B",
		4053 =>	x"0B000000",
		4054 =>	x"00000000",
		4055 =>	x"0C0C0D0D",
		4056 =>	x"0C0B0B0B",
		4057 =>	x"0B0D0D00",
		4058 =>	x"00000000",
		4059 =>	x"00000C0C",
		4060 =>	x"0C0C0B0B",
		4061 =>	x"0B000000",
		4062 =>	x"00000000",
		4063 =>	x"0C0C0D0D",
		4064 =>	x"0C0B0B0B",
		4065 =>	x"0B0D0D00",
		4066 =>	x"00000000",
		4067 =>	x"00000D0D",
		4068 =>	x"0C0B0B0B",
		4069 =>	x"0B000000",
		4070 =>	x"00000000",
		4071 =>	x"00000C0C",
		4072 =>	x"000C0C0C",
		4073 =>	x"0C0C0000",
		4074 =>	x"00000000",
		4075 =>	x"00000C00",
		4076 =>	x"00000C0C",
		4077 =>	x"0C0C0C0C",
		4078 =>	x"0C0C0C00",
		4079 =>	x"00000000",
		4080 =>	x"00000C0C",
		4081 =>	x"0C0D0D0C",
		4082 =>	x"0D0D0C0C",
		4083 =>	x"00000000",
		4084 =>	x"0000000C",
		4085 =>	x"0C0C0C0D",
		4086 =>	x"0D0D0C0C",
		4087 =>	x"00000000",
		4088 =>	x"0000000C",
		4089 =>	x"00000C0C",
		4090 =>	x"0C0C0C00",
		4091 =>	x"00000000",
		4092 =>	x"00000000",
		4093 =>	x"00000000",
		4094 =>	x"00000000",
		4095 =>	x"00000000", -- IMG_16x16_muva_pola10
		4096 =>	x"00000000",
		4097 =>	x"000C0000",
		4098 =>	x"00000000",
		4099 =>	x"0000000C",
		4100 =>	x"00000000",
		4101 =>	x"0C0C0C00",
		4102 =>	x"00000000",
		4103 =>	x"0000000C",
		4104 =>	x"0C000C0C",
		4105 =>	x"0C0C0C0C",
		4106 =>	x"0C000000",
		4107 =>	x"0000000D",
		4108 =>	x"0C000C0C",
		4109 =>	x"0C0C0C0C",
		4110 =>	x"0C000000",
		4111 =>	x"00000C0D",
		4112 =>	x"0D0C0B0B",
		4113 =>	x"0C000000",
		4114 =>	x"0C0C0000",
		4115 =>	x"00000C0C",
		4116 =>	x"0C0B0B0B",
		4117 =>	x"0B0B0000",
		4118 =>	x"0C0C0C00",
		4119 =>	x"000C0D0D",
		4120 =>	x"0C0C0B0B",
		4121 =>	x"0B0D0D00",
		4122 =>	x"000C0C00",
		4123 =>	x"00000D0D",
		4124 =>	x"0C0B0B0B",
		4125 =>	x"0B000000",
		4126 =>	x"00000C0C",
		4127 =>	x"00000C00",
		4128 =>	x"0C0B0B0B",
		4129 =>	x"0B0D0D00",
		4130 =>	x"00000000",
		4131 =>	x"000C0000",
		4132 =>	x"0C0C0C0B",
		4133 =>	x"00000000",
		4134 =>	x"00000C00",
		4135 =>	x"00000000",
		4136 =>	x"0C0C0C00",
		4137 =>	x"00000C00",
		4138 =>	x"0C0C0000",
		4139 =>	x"00000000",
		4140 =>	x"000C0C0C",
		4141 =>	x"0C0C0C0C",
		4142 =>	x"0C000000",
		4143 =>	x"00000000",
		4144 =>	x"00000C0C",
		4145 =>	x"0C0C0C0C",
		4146 =>	x"00000000",
		4147 =>	x"00000000",
		4148 =>	x"000C0000",
		4149 =>	x"00000000",
		4150 =>	x"00000000",
		4151 =>	x"00000000",
		4152 =>	x"00000000",
		4153 =>	x"00000000",
		4154 =>	x"00000000",
		4155 =>	x"00000000",
		4156 =>	x"00000000",
		4157 =>	x"00000000",
		4158 =>	x"00000000",
		4159 =>	x"00000000", -- IMG_16x16_muva_pola11
		4160 =>	x"0000000C",
		4161 =>	x"00000000",
		4162 =>	x"00000000",
		4163 =>	x"00000000",
		4164 =>	x"0000000C",
		4165 =>	x"00000000",
		4166 =>	x"00000000",
		4167 =>	x"00000000",
		4168 =>	x"0C0D0D00",
		4169 =>	x"000C0C00",
		4170 =>	x"0C0C0000",
		4171 =>	x"0000000C",
		4172 =>	x"000D0D0C",
		4173 =>	x"0C0C0C0C",
		4174 =>	x"0C000000",
		4175 =>	x"0000000D",
		4176 =>	x"0D0C0C0B",
		4177 =>	x"0B0C0C0C",
		4178 =>	x"0C000000",
		4179 =>	x"0000000D",
		4180 =>	x"0D0C0C0B",
		4181 =>	x"0B0B000C",
		4182 =>	x"0C0C0000",
		4183 =>	x"000C0C00",
		4184 =>	x"0C0B0B0B",
		4185 =>	x"0B0B0B00",
		4186 =>	x"0C0C0C00",
		4187 =>	x"00000000",
		4188 =>	x"0C0B0B0B",
		4189 =>	x"0B0B0D00",
		4190 =>	x"0C0C0C00",
		4191 =>	x"0000000C",
		4192 =>	x"0C0C0B0B",
		4193 =>	x"0B000D00",
		4194 =>	x"000C0C00",
		4195 =>	x"0000000C",
		4196 =>	x"0C0C000B",
		4197 =>	x"0D0D0000",
		4198 =>	x"000C0C00",
		4199 =>	x"00000000",
		4200 =>	x"0C0C0C00",
		4201 =>	x"00000000",
		4202 =>	x"000C0000",
		4203 =>	x"0000000C",
		4204 =>	x"0C0C0C0C",
		4205 =>	x"0C000000",
		4206 =>	x"000C0000",
		4207 =>	x"0000000C",
		4208 =>	x"00000C0C",
		4209 =>	x"0C0C0C0C",
		4210 =>	x"0C000000",
		4211 =>	x"00000000",
		4212 =>	x"0000000C",
		4213 =>	x"0C0C0C00",
		4214 =>	x"00000000",
		4215 =>	x"00000000",
		4216 =>	x"00000000",
		4217 =>	x"00000000",
		4218 =>	x"00000000",
		4219 =>	x"00000000",
		4220 =>	x"00000000",
		4221 =>	x"00000000",
		4222 =>	x"00000000",
		4223 =>	x"00000000", -- IMG_16x16_muva_pola12
		4224 =>	x"0000000C",
		4225 =>	x"00000C00",
		4226 =>	x"00000000",
		4227 =>	x"00000000",
		4228 =>	x"000C0C0D",
		4229 =>	x"0D0C0000",
		4230 =>	x"00000000",
		4231 =>	x"00000C0C",
		4232 =>	x"0D0D0C0D",
		4233 =>	x"0D000000",
		4234 =>	x"00000000",
		4235 =>	x"0000000C",
		4236 =>	x"0C0D0C0C",
		4237 =>	x"0C0C0C0C",
		4238 =>	x"00000000",
		4239 =>	x"00000000",
		4240 =>	x"000C0B0C",
		4241 =>	x"0B0B0C0C",
		4242 =>	x"0C000C00",
		4243 =>	x"0000000C",
		4244 =>	x"0C0B0B0B",
		4245 =>	x"0B0B0C0C",
		4246 =>	x"0C0C0000",
		4247 =>	x"0000000C",
		4248 =>	x"0C0B0B0B",
		4249 =>	x"0B0B0B00",
		4250 =>	x"0C0C0000",
		4251 =>	x"00000C0C",
		4252 =>	x"0C0C0B0B",
		4253 =>	x"0B0B0000",
		4254 =>	x"0C0C0000",
		4255 =>	x"000C0C0C",
		4256 =>	x"0C000B0D",
		4257 =>	x"000D0000",
		4258 =>	x"0C0C0000",
		4259 =>	x"00000C0C",
		4260 =>	x"0C00000D",
		4261 =>	x"000D000C",
		4262 =>	x"0C0C0000",
		4263 =>	x"0000000C",
		4264 =>	x"0C000000",
		4265 =>	x"00000000",
		4266 =>	x"0C0C0000",
		4267 =>	x"0000000C",
		4268 =>	x"0C0C0C00",
		4269 =>	x"0000000C",
		4270 =>	x"0C000000",
		4271 =>	x"00000000",
		4272 =>	x"000C0C0C",
		4273 =>	x"0000000C",
		4274 =>	x"00000000",
		4275 =>	x"00000000",
		4276 =>	x"00000C0C",
		4277 =>	x"0C000C00",
		4278 =>	x"00000000",
		4279 =>	x"00000000",
		4280 =>	x"00000000",
		4281 =>	x"0C000000",
		4282 =>	x"00000000",
		4283 =>	x"00000000",
		4284 =>	x"00000000",
		4285 =>	x"00000000",
		4286 =>	x"00000000",


--			***** MAP *****


		4287 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4288 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4289 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4290 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4291 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4292 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4293 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4294 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4295 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4296 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4297 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4298 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4299 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4300 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4301 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4302 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4303 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4304 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4305 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4306 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4307 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4308 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4309 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4310 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4311 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4312 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4313 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4314 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4315 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4316 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4317 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4318 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4319 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4320 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4321 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4322 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4323 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4324 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4325 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4326 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4327 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4328 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4329 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4330 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4331 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4332 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4333 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4334 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4335 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4336 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4337 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4338 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4339 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4340 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4341 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4342 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4343 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4344 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4345 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4346 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4347 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4348 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4349 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4350 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4351 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4352 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4353 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4354 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4355 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4356 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4357 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4358 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4359 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4360 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4361 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4362 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4363 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4364 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4365 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4366 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4367 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4368 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4369 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4370 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4371 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4372 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4373 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4374 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4375 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4376 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4377 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4378 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4379 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4380 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4381 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4382 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4383 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4384 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4385 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4386 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4387 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4388 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4389 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4390 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4391 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4392 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4393 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4394 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4395 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4396 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4397 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4398 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4399 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4400 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4401 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4402 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4403 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4404 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4405 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4406 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4407 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4408 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4409 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4410 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4411 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4412 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4413 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4414 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4415 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4416 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4417 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4418 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4419 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4420 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4421 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4422 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4423 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4424 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4425 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4426 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4427 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4428 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4429 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4430 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4431 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4432 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4433 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4434 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4435 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4436 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4437 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4438 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4439 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4440 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4441 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4442 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4443 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4444 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4445 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4446 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4447 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4448 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4449 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4450 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4451 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4452 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4453 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4454 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4455 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4456 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4457 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4458 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4459 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4460 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4461 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4462 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4463 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4464 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4465 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4466 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4467 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4468 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4469 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4470 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4471 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4472 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4473 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4474 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4475 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4476 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4477 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4478 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4479 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4480 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4481 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4482 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4483 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4484 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4485 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4486 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4487 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4488 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4489 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4490 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4491 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4492 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4493 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4494 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4495 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4496 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4497 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4498 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4499 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4500 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4501 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4502 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4503 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4504 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4505 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4506 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4507 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4508 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4509 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4510 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4511 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4512 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4513 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4514 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4515 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4516 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4517 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4518 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4519 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4520 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4521 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4522 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4523 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4524 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4525 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4526 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4527 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4528 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4529 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4530 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4531 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4532 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4533 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4534 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4535 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4536 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4537 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4538 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4539 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4540 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4541 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4542 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4543 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4544 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4545 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4546 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4547 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4548 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4549 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4550 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4551 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4552 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4553 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4554 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4555 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4556 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4557 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4558 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4559 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4560 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4561 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4562 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4563 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4564 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4565 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4566 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4567 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4568 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4569 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4570 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4571 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4572 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4573 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4574 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4575 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4576 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4577 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4578 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4579 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4580 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4581 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4582 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4583 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4584 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4585 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4586 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4587 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4588 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4589 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4590 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4591 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4592 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4593 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4594 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4595 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4596 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4597 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4598 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4599 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4600 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4601 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4602 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4603 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4604 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4605 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4606 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4607 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4608 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4609 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4610 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4611 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4612 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4613 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4614 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4615 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4616 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4617 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4618 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4619 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4620 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4621 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4622 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4623 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4624 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4625 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4626 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4627 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4628 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4629 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4630 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4631 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4632 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4633 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4634 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4635 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4636 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4637 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4638 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4639 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4640 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4641 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4642 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4643 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4644 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4645 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4646 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4647 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4648 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4649 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4650 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4651 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4652 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4653 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4654 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4655 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4656 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4657 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4658 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4659 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4660 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4661 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4662 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4663 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4664 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4665 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4666 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4667 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4668 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4669 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4670 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4671 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4672 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4673 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4674 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4675 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4676 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4677 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4678 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4679 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4680 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4681 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4682 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4683 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4684 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4685 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4686 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4687 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4688 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4689 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4690 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4691 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4692 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4693 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4694 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4695 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4696 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4697 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4698 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4699 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4700 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4701 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4702 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4703 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4704 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4705 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4706 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4707 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4708 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4709 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4710 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4711 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4712 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4713 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4714 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4715 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4716 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4717 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4718 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4719 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4720 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4721 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4722 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4723 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4724 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4725 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4726 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4727 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4728 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4729 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4730 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4731 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4732 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4733 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4734 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4735 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4736 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4737 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4738 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4739 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4740 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4741 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4742 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4743 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4744 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4745 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4746 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4747 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4748 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4749 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4750 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4751 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4752 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4753 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4754 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4755 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4756 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4757 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4758 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4759 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4760 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4761 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4762 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4763 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4764 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4765 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4766 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4767 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4768 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4769 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4770 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4771 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4772 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4773 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4774 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4775 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4776 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4777 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4778 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4779 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4780 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4781 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4782 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4783 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4784 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4785 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4786 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4787 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4788 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4789 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4790 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4791 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4792 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4793 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4794 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4795 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4796 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4797 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4798 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4799 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4800 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4801 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4802 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4803 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4804 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4805 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4806 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4807 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4808 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4809 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4810 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4811 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4812 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4813 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4814 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4815 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4816 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4817 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4818 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4819 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4820 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4821 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4822 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4823 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4824 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4825 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4826 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4827 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4828 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4829 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4830 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4831 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4832 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4833 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4834 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4835 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4836 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4837 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4838 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4839 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4840 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4841 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4842 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4843 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4844 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4845 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4846 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4847 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4848 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4849 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4850 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4851 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4852 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4853 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4854 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4855 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4856 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4857 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4858 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4859 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4860 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4861 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4862 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4863 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4864 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4865 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4866 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4867 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4868 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4869 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4870 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4871 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4872 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4873 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4874 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4875 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4876 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4877 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4878 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4879 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4880 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4881 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4882 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4883 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4884 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4885 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4886 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4887 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4888 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4889 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4890 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4891 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4892 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4893 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4894 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4895 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4896 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4897 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4898 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4899 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4900 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4901 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4902 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4903 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4904 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4905 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4906 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4907 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4908 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4909 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4910 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4911 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4912 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4913 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4914 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4915 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4916 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4917 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4918 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4919 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4920 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4921 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4922 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4923 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4924 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4925 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4926 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4927 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4928 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4929 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4930 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4931 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4932 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4933 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4934 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4935 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4936 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4937 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4938 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4939 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4940 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4941 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4942 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4943 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4944 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4945 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4946 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4947 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4948 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4949 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4950 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4951 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4952 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4953 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4954 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4955 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4956 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4957 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4958 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4959 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4960 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4961 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4962 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4963 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4964 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4965 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4966 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4967 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4968 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4969 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4970 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4971 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4972 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4973 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4974 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4975 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4976 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4977 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4978 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4979 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4980 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4981 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4982 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4983 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4984 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4985 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4986 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4987 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4988 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4989 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4990 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4991 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4992 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4993 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4994 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4995 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4996 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4997 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4998 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		4999 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5000 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5001 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5002 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5003 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5004 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5005 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5006 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5007 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5008 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5009 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5010 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5011 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5012 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5013 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5014 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5015 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5016 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5017 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5018 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5019 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5020 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5021 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5022 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5023 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5024 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5025 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5026 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5027 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5028 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5029 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5030 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5031 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5032 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5033 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5034 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5035 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5036 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5037 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5038 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5039 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5040 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5041 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5042 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5043 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5044 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5045 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5046 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5047 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5048 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5049 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5050 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5051 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5052 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5053 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5054 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5055 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5056 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5057 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5058 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5059 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5060 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5061 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5062 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5063 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5064 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5065 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5066 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5067 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5068 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5069 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5070 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5071 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5072 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5073 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5074 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5075 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5076 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5077 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5078 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5079 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5080 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5081 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5082 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5083 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5084 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5085 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5086 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5087 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5088 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5089 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5090 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5091 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5092 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5093 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5094 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5095 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5096 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5097 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5098 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5099 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5100 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5101 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5102 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5103 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5104 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5105 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5106 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5107 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5108 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5109 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5110 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5111 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5112 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5113 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5114 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5115 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5116 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5117 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5118 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5119 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5120 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5121 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5122 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5123 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5124 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5125 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5126 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5127 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5128 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5129 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5130 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5131 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5132 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5133 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5134 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5135 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5136 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5137 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5138 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5139 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5140 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5141 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5142 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5143 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5144 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5145 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5146 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5147 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5148 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5149 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5150 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5151 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5152 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5153 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5154 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5155 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5156 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5157 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5158 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5159 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5160 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5161 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5162 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5163 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5164 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5165 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5166 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5167 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5168 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5169 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5170 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5171 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5172 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5173 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5174 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5175 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5176 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5177 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5178 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5179 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5180 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5181 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5182 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5183 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5184 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5185 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5186 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5187 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5188 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5189 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5190 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5191 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5192 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5193 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5194 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5195 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5196 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5197 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5198 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5199 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5200 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5201 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5202 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5203 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5204 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5205 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5206 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5207 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5208 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5209 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5210 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5211 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5212 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5213 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5214 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5215 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5216 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5217 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5218 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5219 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5220 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5221 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5222 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5223 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5224 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5225 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5226 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5227 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5228 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5229 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5230 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5231 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5232 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5233 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5234 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5235 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5236 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5237 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5238 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5239 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5240 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5241 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5242 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5243 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5244 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5245 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5246 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5247 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5248 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5249 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5250 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5251 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5252 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5253 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5254 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5255 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5256 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5257 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5258 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5259 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5260 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5261 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5262 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5263 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5264 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5265 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5266 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5267 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5268 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5269 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5270 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5271 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5272 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5273 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5274 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5275 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5276 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5277 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5278 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5279 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5280 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5281 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5282 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5283 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5284 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5285 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5286 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5287 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5288 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5289 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5290 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5291 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5292 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5293 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5294 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5295 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5296 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5297 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5298 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5299 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5300 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5301 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5302 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5303 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5304 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5305 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5306 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5307 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5308 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5309 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5310 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5311 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5312 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5313 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5314 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5315 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5316 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5317 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5318 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5319 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5320 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5321 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5322 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5323 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5324 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5325 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5326 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5327 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5328 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5329 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5330 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5331 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5332 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5333 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5334 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5335 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5336 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5337 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5338 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5339 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5340 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5341 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5342 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5343 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5344 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5345 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5346 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5347 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5348 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5349 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5350 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5351 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5352 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5353 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5354 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5355 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5356 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5357 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5358 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5359 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5360 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5361 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5362 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5363 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5364 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5365 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5366 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5367 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5368 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5369 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5370 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5371 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5372 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5373 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5374 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5375 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5376 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5377 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5378 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5379 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5380 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5381 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5382 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5383 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5384 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5385 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5386 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5387 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5388 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5389 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5390 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5391 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5392 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5393 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5394 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5395 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5396 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5397 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5398 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5399 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5400 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5401 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5402 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5403 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5404 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5405 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5406 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5407 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5408 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5409 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5410 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5411 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5412 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5413 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5414 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5415 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5416 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5417 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5418 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5419 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5420 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5421 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5422 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5423 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5424 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5425 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5426 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5427 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5428 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5429 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5430 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5431 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5432 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5433 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5434 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5435 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5436 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5437 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5438 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5439 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5440 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5441 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5442 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5443 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5444 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5445 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5446 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5447 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5448 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5449 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5450 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5451 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5452 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5453 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5454 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5455 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5456 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5457 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5458 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5459 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5460 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5461 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5462 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5463 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5464 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5465 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5466 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5467 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5468 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5469 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5470 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5471 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5472 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5473 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5474 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5475 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5476 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5477 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5478 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5479 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5480 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5481 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5482 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5483 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5484 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5485 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5486 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5487 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5488 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5489 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5490 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5491 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5492 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5493 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5494 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5495 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5496 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5497 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5498 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5499 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5500 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5501 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5502 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5503 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5504 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5505 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5506 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5507 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5508 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5509 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5510 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5511 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5512 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5513 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5514 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5515 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5516 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5517 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5518 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5519 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5520 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5521 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5522 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5523 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5524 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5525 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5526 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5527 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5528 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5529 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5530 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5531 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5532 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5533 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5534 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5535 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5536 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5537 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5538 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5539 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5540 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5541 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5542 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5543 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5544 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5545 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5546 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5547 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5548 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5549 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5550 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5551 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5552 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5553 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5554 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5555 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5556 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5557 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5558 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5559 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5560 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5561 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5562 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5563 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5564 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5565 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5566 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5567 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5568 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5569 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5570 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5571 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5572 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5573 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5574 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5575 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5576 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5577 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5578 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5579 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5580 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5581 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5582 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5583 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5584 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5585 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5586 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5587 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5588 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5589 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5590 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5591 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5592 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5593 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5594 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5595 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5596 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5597 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5598 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5599 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5600 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5601 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5602 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5603 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5604 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5605 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5606 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5607 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5608 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5609 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5610 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5611 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5612 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5613 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5614 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5615 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5616 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5617 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5618 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5619 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5620 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5621 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5622 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5623 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5624 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5625 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5626 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5627 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5628 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5629 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5630 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5631 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5632 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5633 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5634 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5635 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5636 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5637 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5638 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5639 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5640 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5641 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5642 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5643 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5644 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5645 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5646 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5647 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5648 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5649 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5650 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5651 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5652 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5653 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5654 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5655 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5656 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5657 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5658 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5659 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5660 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5661 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5662 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5663 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5664 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5665 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5666 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5667 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5668 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5669 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5670 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5671 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5672 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5673 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5674 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5675 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5676 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5677 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5678 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5679 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5680 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5681 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5682 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5683 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5684 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5685 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5686 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5687 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5688 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5689 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5690 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5691 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5692 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5693 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5694 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5695 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5696 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5697 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5698 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5699 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5700 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5701 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5702 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5703 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5704 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5705 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5706 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5707 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5708 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5709 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5710 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5711 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5712 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5713 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5714 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5715 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5716 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5717 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5718 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5719 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5720 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5721 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5722 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5723 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5724 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5725 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5726 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5727 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5728 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5729 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5730 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5731 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5732 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5733 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5734 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5735 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5736 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5737 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5738 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5739 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5740 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5741 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5742 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5743 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5744 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5745 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5746 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5747 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5748 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5749 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5750 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5751 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5752 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5753 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5754 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5755 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5756 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5757 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5758 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5759 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5760 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5761 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5762 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5763 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5764 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5765 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5766 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5767 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5768 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5769 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5770 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5771 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5772 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5773 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5774 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5775 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5776 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5777 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5778 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5779 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5780 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5781 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5782 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5783 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5784 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5785 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5786 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5787 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5788 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5789 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5790 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5791 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5792 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5793 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5794 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5795 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5796 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5797 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5798 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5799 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5800 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5801 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5802 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5803 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5804 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5805 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5806 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5807 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5808 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5809 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5810 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5811 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5812 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5813 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5814 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5815 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5816 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5817 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5818 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5819 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5820 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5821 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5822 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5823 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5824 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5825 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5826 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5827 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5828 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5829 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5830 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5831 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5832 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5833 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5834 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5835 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5836 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5837 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5838 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5839 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5840 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5841 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5842 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5843 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5844 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5845 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5846 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5847 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5848 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5849 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5850 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5851 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5852 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5853 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5854 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5855 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5856 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5857 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5858 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5859 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5860 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5861 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5862 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5863 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5864 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5865 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5866 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5867 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5868 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5869 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5870 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5871 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5872 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5873 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5874 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5875 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5876 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5877 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5878 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5879 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5880 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5881 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5882 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5883 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5884 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5885 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5886 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5887 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5888 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5889 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5890 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5891 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5892 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5893 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5894 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5895 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5896 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5897 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5898 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5899 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5900 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5901 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5902 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5903 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5904 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5905 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5906 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5907 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5908 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5909 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5910 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5911 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5912 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5913 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5914 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5915 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5916 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5917 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5918 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5919 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5920 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5921 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5922 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5923 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5924 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5925 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5926 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5927 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5928 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5929 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5930 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5931 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5932 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5933 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5934 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5935 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5936 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5937 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5938 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5939 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5940 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5941 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5942 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5943 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5944 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5945 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5946 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5947 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5948 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5949 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5950 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5951 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5952 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5953 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5954 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5955 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5956 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5957 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5958 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5959 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5960 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5961 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5962 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5963 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5964 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5965 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5966 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5967 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5968 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5969 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5970 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5971 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5972 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5973 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5974 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5975 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5976 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5977 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5978 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5979 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5980 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5981 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5982 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5983 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5984 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5985 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5986 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5987 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5988 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5989 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5990 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5991 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5992 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5993 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5994 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5995 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5996 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5997 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5998 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		5999 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6000 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6001 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6002 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6003 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6004 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6005 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6006 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6007 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6008 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6009 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6010 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6011 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6012 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6013 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6014 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6015 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6016 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6017 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6018 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6019 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6020 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6021 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6022 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6023 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6024 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6025 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6026 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6027 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6028 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6029 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6030 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6031 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6032 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6033 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6034 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6035 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6036 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6037 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6038 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6039 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6040 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6041 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6042 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6043 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6044 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6045 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6046 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6047 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6048 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6049 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6050 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6051 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6052 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6053 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6054 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6055 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6056 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6057 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6058 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6059 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6060 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6061 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6062 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6063 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6064 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6065 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6066 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6067 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6068 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6069 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6070 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6071 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6072 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6073 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6074 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6075 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6076 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6077 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6078 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6079 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6080 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6081 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6082 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6083 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6084 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6085 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6086 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6087 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6088 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6089 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6090 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6091 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6092 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6093 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6094 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6095 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6096 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6097 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6098 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6099 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6100 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6101 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6102 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6103 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6104 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6105 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6106 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6107 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6108 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6109 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6110 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6111 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6112 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6113 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6114 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6115 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6116 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6117 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6118 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6119 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6120 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6121 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6122 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6123 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6124 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6125 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6126 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6127 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6128 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6129 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6130 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6131 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6132 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6133 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6134 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6135 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6136 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6137 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6138 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6139 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6140 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6141 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6142 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6143 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6144 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6145 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6146 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6147 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6148 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6149 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6150 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6151 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6152 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6153 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6154 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6155 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6156 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6157 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6158 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6159 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6160 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6161 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6162 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6163 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6164 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6165 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6166 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6167 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6168 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6169 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6170 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6171 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6172 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6173 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6174 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6175 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6176 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6177 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6178 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6179 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6180 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6181 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6182 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6183 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6184 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6185 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6186 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6187 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6188 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6189 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6190 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6191 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6192 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6193 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6194 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6195 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6196 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6197 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6198 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6199 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6200 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6201 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6202 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6203 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6204 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6205 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6206 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6207 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6208 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6209 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6210 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6211 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6212 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6213 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6214 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6215 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6216 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6217 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6218 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6219 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6220 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6221 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6222 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6223 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6224 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6225 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6226 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6227 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6228 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6229 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6230 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6231 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6232 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6233 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6234 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6235 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6236 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6237 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6238 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6239 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6240 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6241 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6242 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6243 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6244 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6245 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6246 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6247 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6248 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6249 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6250 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6251 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6252 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6253 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6254 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6255 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6256 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6257 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6258 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6259 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6260 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6261 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6262 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6263 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6264 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6265 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6266 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6267 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6268 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6269 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6270 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6271 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6272 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6273 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6274 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6275 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6276 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6277 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6278 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6279 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6280 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6281 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6282 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6283 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6284 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6285 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6286 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6287 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6288 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6289 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6290 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6291 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6292 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6293 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6294 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6295 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6296 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6297 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6298 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6299 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6300 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6301 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6302 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6303 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6304 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6305 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6306 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6307 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6308 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6309 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6310 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6311 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6312 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6313 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6314 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6315 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6316 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6317 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6318 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6319 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6320 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6321 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6322 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6323 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6324 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6325 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6326 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6327 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6328 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6329 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6330 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6331 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6332 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6333 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6334 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6335 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6336 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6337 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6338 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6339 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6340 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6341 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6342 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6343 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6344 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6345 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6346 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6347 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6348 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6349 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6350 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6351 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6352 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6353 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6354 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6355 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6356 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6357 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6358 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6359 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6360 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6361 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6362 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6363 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6364 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6365 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6366 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6367 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6368 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6369 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6370 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6371 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6372 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6373 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6374 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6375 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6376 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6377 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6378 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6379 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6380 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6381 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6382 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6383 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6384 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6385 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6386 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6387 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6388 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6389 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6390 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6391 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6392 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6393 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6394 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6395 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6396 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6397 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6398 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6399 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6400 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6401 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6402 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6403 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6404 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6405 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6406 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6407 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6408 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6409 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6410 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6411 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6412 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6413 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6414 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6415 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6416 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6417 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6418 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6419 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6420 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6421 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6422 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6423 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6424 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6425 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6426 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6427 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6428 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6429 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6430 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6431 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6432 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6433 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6434 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6435 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6436 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6437 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6438 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6439 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6440 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6441 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6442 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6443 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6444 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6445 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6446 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6447 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6448 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6449 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6450 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6451 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6452 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6453 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6454 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6455 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6456 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6457 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6458 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6459 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6460 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6461 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6462 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6463 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6464 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6465 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6466 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6467 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6468 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6469 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6470 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6471 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6472 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6473 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6474 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6475 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6476 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6477 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6478 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6479 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6480 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6481 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6482 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6483 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6484 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6485 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6486 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6487 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6488 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6489 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6490 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6491 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6492 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6493 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6494 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6495 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6496 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6497 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6498 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6499 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6500 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6501 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6502 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6503 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6504 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6505 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6506 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6507 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6508 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6509 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6510 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6511 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6512 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6513 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6514 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6515 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6516 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6517 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6518 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6519 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6520 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6521 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6522 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6523 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6524 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6525 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6526 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6527 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6528 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6529 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6530 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6531 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6532 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6533 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6534 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6535 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6536 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6537 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6538 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6539 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6540 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6541 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6542 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6543 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6544 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6545 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6546 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6547 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6548 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6549 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6550 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6551 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6552 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6553 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6554 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6555 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6556 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6557 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6558 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6559 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6560 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6561 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6562 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6563 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6564 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6565 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6566 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6567 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6568 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6569 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6570 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6571 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6572 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6573 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6574 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6575 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6576 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6577 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6578 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6579 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6580 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6581 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6582 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6583 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6584 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6585 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6586 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6587 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6588 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6589 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6590 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6591 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6592 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6593 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6594 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6595 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6596 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6597 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6598 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6599 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6600 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6601 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6602 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6603 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6604 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6605 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6606 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6607 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6608 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6609 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6610 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6611 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6612 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6613 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6614 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6615 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6616 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6617 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6618 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6619 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6620 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6621 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6622 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6623 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6624 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6625 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6626 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6627 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6628 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6629 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6630 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6631 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6632 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6633 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6634 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6635 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6636 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6637 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6638 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6639 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6640 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6641 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6642 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6643 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6644 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6645 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6646 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6647 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6648 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6649 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6650 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6651 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6652 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6653 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6654 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6655 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6656 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6657 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6658 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6659 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6660 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6661 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6662 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6663 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6664 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6665 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6666 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6667 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6668 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6669 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6670 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6671 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6672 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6673 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6674 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6675 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6676 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6677 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6678 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6679 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6680 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6681 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6682 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6683 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6684 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6685 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6686 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6687 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6688 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6689 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6690 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6691 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6692 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6693 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6694 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6695 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6696 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6697 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6698 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6699 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6700 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6701 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6702 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6703 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6704 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6705 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6706 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6707 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6708 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6709 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6710 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6711 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6712 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6713 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6714 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6715 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6716 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6717 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6718 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6719 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6720 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6721 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6722 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6723 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6724 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6725 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6726 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6727 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6728 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6729 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6730 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6731 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6732 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6733 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6734 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6735 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6736 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6737 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6738 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6739 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6740 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6741 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6742 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6743 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6744 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6745 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6746 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6747 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6748 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6749 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6750 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6751 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6752 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6753 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6754 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6755 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6756 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6757 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6758 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6759 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6760 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6761 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6762 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6763 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6764 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6765 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6766 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6767 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6768 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6769 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6770 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6771 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6772 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6773 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6774 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6775 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6776 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6777 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6778 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6779 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6780 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6781 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6782 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6783 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6784 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6785 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6786 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6787 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6788 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6789 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6790 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6791 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6792 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6793 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6794 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6795 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6796 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6797 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6798 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6799 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6800 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6801 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6802 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6803 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6804 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6805 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6806 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6807 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6808 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6809 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6810 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6811 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6812 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6813 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6814 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6815 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6816 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6817 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6818 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6819 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6820 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6821 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6822 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6823 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6824 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6825 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6826 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6827 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6828 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6829 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6830 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6831 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6832 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6833 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6834 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6835 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6836 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6837 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6838 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6839 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6840 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6841 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6842 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6843 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6844 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6845 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6846 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6847 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6848 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6849 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6850 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6851 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6852 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6853 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6854 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6855 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6856 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6857 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6858 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6859 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6860 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6861 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6862 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6863 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6864 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6865 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6866 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6867 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6868 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6869 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6870 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6871 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6872 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6873 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6874 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6875 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6876 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6877 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6878 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6879 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6880 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6881 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6882 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6883 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6884 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6885 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6886 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6887 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6888 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6889 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6890 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6891 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6892 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6893 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6894 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6895 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6896 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6897 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6898 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6899 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6900 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6901 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6902 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6903 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6904 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6905 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6906 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6907 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6908 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6909 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6910 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6911 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6912 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6913 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6914 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6915 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6916 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6917 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6918 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6919 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6920 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6921 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6922 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6923 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6924 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6925 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6926 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6927 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6928 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6929 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6930 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6931 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6932 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6933 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6934 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6935 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6936 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6937 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6938 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6939 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6940 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6941 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6942 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6943 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6944 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6945 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6946 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6947 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6948 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6949 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6950 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6951 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6952 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6953 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6954 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6955 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6956 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6957 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6958 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6959 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6960 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6961 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6962 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6963 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6964 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6965 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6966 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6967 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6968 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6969 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6970 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6971 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6972 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6973 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6974 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6975 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6976 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6977 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6978 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6979 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6980 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6981 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6982 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6983 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6984 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6985 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6986 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6987 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6988 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6989 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6990 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6991 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6992 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6993 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6994 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6995 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6996 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6997 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6998 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		6999 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7000 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7001 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7002 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7003 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7004 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7005 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7006 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7007 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7008 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7009 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7010 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7011 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7012 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7013 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7014 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7015 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7016 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7017 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7018 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7019 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7020 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7021 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7022 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7023 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7024 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7025 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7026 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7027 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7028 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7029 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7030 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7031 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7032 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7033 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7034 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7035 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7036 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7037 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7038 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7039 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7040 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7041 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7042 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7043 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7044 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7045 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7046 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7047 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7048 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7049 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7050 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7051 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7052 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7053 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7054 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7055 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7056 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7057 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7058 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7059 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7060 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7061 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7062 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7063 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7064 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7065 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7066 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7067 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7068 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7069 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7070 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7071 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7072 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7073 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7074 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7075 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7076 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7077 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7078 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7079 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7080 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7081 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7082 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7083 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7084 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7085 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7086 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7087 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7088 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7089 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7090 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7091 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7092 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7093 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7094 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7095 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7096 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7097 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7098 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7099 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7100 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7101 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7102 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7103 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7104 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7105 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7106 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7107 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7108 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7109 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7110 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7111 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7112 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7113 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7114 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7115 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7116 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7117 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7118 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7119 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7120 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7121 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7122 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7123 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7124 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7125 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7126 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7127 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7128 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7129 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7130 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7131 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7132 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7133 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7134 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7135 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7136 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7137 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7138 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7139 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7140 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7141 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7142 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7143 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7144 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7145 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7146 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7147 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7148 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7149 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7150 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7151 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7152 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7153 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7154 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7155 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7156 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7157 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7158 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7159 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7160 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7161 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7162 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7163 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7164 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7165 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7166 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7167 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7168 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7169 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7170 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7171 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7172 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7173 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7174 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7175 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7176 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7177 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7178 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7179 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7180 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7181 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7182 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7183 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7184 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7185 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7186 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7187 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7188 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7189 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7190 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7191 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7192 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7193 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7194 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7195 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7196 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7197 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7198 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7199 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7200 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7201 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7202 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7203 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7204 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7205 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7206 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7207 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7208 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7209 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7210 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7211 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7212 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7213 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7214 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7215 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7216 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7217 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7218 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7219 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7220 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7221 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7222 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7223 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7224 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7225 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7226 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7227 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7228 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7229 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7230 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7231 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7232 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7233 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7234 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7235 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7236 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7237 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7238 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7239 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7240 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7241 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7242 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7243 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7244 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7245 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7246 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7247 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7248 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7249 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7250 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7251 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7252 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7253 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7254 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7255 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7256 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7257 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7258 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7259 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7260 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7261 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7262 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7263 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7264 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7265 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7266 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7267 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7268 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7269 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7270 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7271 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7272 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7273 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7274 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7275 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7276 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7277 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7278 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7279 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7280 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7281 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7282 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7283 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7284 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7285 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7286 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7287 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7288 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7289 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7290 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7291 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7292 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7293 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7294 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7295 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7296 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7297 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7298 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7299 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7300 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7301 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7302 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7303 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7304 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7305 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7306 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7307 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7308 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7309 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7310 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7311 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7312 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7313 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7314 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7315 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7316 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7317 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7318 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7319 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7320 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7321 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7322 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7323 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7324 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7325 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7326 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7327 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7328 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7329 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7330 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7331 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7332 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7333 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7334 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7335 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7336 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7337 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7338 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7339 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7340 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7341 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7342 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7343 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7344 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7345 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7346 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7347 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7348 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7349 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7350 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7351 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7352 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7353 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7354 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7355 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7356 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7357 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7358 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7359 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7360 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7361 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7362 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7363 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7364 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7365 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7366 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7367 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7368 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7369 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7370 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7371 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7372 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7373 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7374 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7375 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7376 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7377 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7378 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7379 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7380 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7381 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7382 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7383 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7384 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7385 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7386 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7387 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7388 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7389 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7390 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7391 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7392 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7393 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7394 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7395 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7396 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7397 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7398 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7399 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7400 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7401 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7402 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7403 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7404 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7405 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7406 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7407 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7408 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7409 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7410 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7411 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7412 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7413 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7414 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7415 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7416 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7417 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7418 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7419 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7420 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7421 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7422 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7423 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7424 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7425 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7426 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7427 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7428 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7429 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7430 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7431 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7432 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7433 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7434 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7435 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7436 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7437 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7438 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7439 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7440 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7441 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7442 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7443 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7444 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7445 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7446 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7447 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7448 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7449 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7450 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7451 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7452 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7453 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7454 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7455 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7456 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7457 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7458 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7459 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7460 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7461 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7462 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7463 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7464 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7465 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7466 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7467 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7468 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7469 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7470 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7471 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7472 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7473 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7474 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7475 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7476 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7477 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7478 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7479 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7480 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7481 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7482 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7483 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7484 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7485 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7486 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7487 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7488 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7489 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7490 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7491 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7492 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7493 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7494 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7495 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7496 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7497 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7498 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7499 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7500 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7501 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7502 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7503 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7504 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7505 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7506 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7507 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7508 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7509 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7510 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7511 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7512 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7513 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7514 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7515 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7516 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7517 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7518 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7519 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7520 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7521 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7522 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7523 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7524 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7525 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7526 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7527 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7528 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7529 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7530 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7531 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7532 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7533 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7534 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7535 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7536 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7537 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7538 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7539 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7540 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7541 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7542 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7543 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7544 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7545 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7546 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7547 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7548 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7549 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7550 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7551 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7552 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7553 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7554 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7555 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7556 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7557 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7558 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7559 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7560 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7561 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7562 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7563 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7564 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7565 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7566 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7567 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7568 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7569 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7570 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7571 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7572 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7573 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7574 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7575 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7576 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7577 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7578 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7579 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7580 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7581 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7582 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7583 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7584 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7585 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7586 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7587 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7588 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7589 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7590 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7591 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7592 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7593 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7594 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7595 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7596 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7597 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7598 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7599 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7600 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7601 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7602 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7603 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7604 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7605 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7606 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7607 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7608 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7609 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7610 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7611 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7612 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7613 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7614 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7615 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7616 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7617 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7618 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7619 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7620 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7621 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7622 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7623 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7624 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7625 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7626 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7627 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7628 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7629 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7630 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7631 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7632 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7633 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7634 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7635 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7636 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7637 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7638 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7639 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7640 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7641 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7642 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7643 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7644 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7645 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7646 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7647 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7648 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7649 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7650 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7651 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7652 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7653 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7654 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7655 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7656 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7657 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7658 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7659 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7660 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7661 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7662 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7663 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7664 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7665 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7666 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7667 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7668 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7669 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7670 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7671 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7672 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7673 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7674 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7675 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7676 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7677 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7678 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7679 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7680 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7681 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7682 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7683 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7684 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7685 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7686 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7687 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7688 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7689 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7690 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7691 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7692 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7693 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7694 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7695 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7696 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7697 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7698 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7699 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7700 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7701 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7702 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7703 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7704 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7705 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7706 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7707 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7708 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7709 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7710 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7711 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7712 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7713 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7714 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7715 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7716 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7717 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7718 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7719 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7720 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7721 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7722 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7723 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7724 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7725 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7726 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7727 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7728 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7729 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7730 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7731 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7732 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7733 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7734 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7735 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7736 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7737 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7738 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7739 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7740 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7741 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7742 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7743 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7744 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7745 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7746 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7747 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7748 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7749 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7750 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7751 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7752 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7753 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7754 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7755 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7756 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7757 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7758 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7759 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7760 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7761 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7762 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7763 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7764 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7765 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7766 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7767 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7768 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7769 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7770 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7771 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7772 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7773 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7774 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7775 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7776 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7777 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7778 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7779 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7780 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7781 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7782 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7783 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7784 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7785 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7786 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7787 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7788 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7789 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7790 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7791 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7792 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7793 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7794 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7795 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7796 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7797 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7798 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7799 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7800 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7801 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7802 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7803 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7804 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7805 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7806 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7807 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7808 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7809 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7810 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7811 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7812 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7813 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7814 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7815 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7816 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7817 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7818 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7819 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7820 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7821 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7822 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7823 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7824 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7825 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7826 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7827 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7828 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7829 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7830 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7831 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7832 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7833 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7834 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7835 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7836 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7837 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7838 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7839 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7840 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7841 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7842 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7843 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7844 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7845 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7846 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7847 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7848 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7849 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7850 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7851 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7852 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7853 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7854 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7855 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7856 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7857 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7858 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7859 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7860 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7861 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7862 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7863 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7864 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7865 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7866 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7867 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7868 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7869 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7870 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7871 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7872 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7873 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7874 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7875 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7876 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7877 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7878 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7879 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7880 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7881 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7882 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7883 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7884 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7885 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7886 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7887 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7888 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7889 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7890 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7891 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7892 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7893 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7894 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7895 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7896 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7897 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7898 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7899 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7900 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7901 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7902 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7903 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7904 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7905 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7906 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7907 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7908 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7909 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7910 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7911 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7912 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7913 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7914 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7915 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7916 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7917 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7918 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7919 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7920 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7921 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7922 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7923 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7924 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7925 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7926 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7927 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7928 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7929 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7930 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7931 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7932 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7933 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7934 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7935 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7936 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7937 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7938 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7939 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7940 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7941 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7942 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7943 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7944 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7945 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7946 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7947 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7948 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7949 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7950 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7951 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7952 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7953 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7954 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7955 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7956 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7957 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7958 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7959 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7960 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7961 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7962 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7963 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7964 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7965 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7966 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7967 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7968 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7969 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7970 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7971 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7972 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7973 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7974 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7975 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7976 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7977 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7978 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7979 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7980 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7981 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7982 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7983 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7984 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7985 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7986 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7987 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7988 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7989 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7990 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7991 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7992 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7993 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7994 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7995 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7996 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7997 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7998 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		7999 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8000 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8001 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8002 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8003 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8004 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8005 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8006 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8007 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8008 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8009 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8010 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8011 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8012 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8013 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8014 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8015 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8016 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8017 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8018 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8019 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8020 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8021 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8022 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8023 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8024 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8025 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8026 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8027 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8028 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8029 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8030 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8031 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8032 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8033 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8034 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8035 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8036 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8037 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8038 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8039 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8040 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8041 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8042 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8043 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8044 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8045 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8046 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8047 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8048 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8049 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8050 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8051 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8052 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8053 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8054 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8055 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8056 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8057 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8058 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8059 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8060 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8061 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8062 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8063 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8064 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8065 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8066 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8067 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8068 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8069 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8070 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8071 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8072 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8073 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8074 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8075 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8076 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8077 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8078 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8079 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8080 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8081 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8082 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8083 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8084 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8085 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8086 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8087 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8088 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8089 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8090 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8091 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8092 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8093 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8094 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8095 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8096 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8097 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8098 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8099 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8100 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8101 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8102 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8103 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8104 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8105 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8106 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8107 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8108 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8109 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8110 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8111 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8112 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8113 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8114 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8115 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8116 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8117 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8118 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8119 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8120 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8121 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8122 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8123 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8124 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8125 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8126 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8127 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8128 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8129 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8130 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8131 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8132 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8133 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8134 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8135 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8136 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8137 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8138 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8139 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8140 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8141 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8142 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8143 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8144 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8145 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8146 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8147 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8148 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8149 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8150 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8151 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8152 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8153 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8154 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8155 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8156 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8157 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8158 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8159 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8160 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8161 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8162 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8163 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8164 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8165 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8166 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8167 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8168 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8169 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8170 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8171 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8172 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8173 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8174 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8175 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8176 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8177 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8178 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8179 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8180 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8181 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8182 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8183 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8184 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8185 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8186 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8187 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8188 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8189 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8190 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8191 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8192 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8193 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8194 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8195 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8196 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8197 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8198 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8199 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8200 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8201 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8202 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8203 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8204 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8205 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8206 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8207 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8208 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8209 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8210 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8211 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8212 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8213 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8214 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8215 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8216 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8217 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8218 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8219 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8220 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8221 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8222 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8223 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8224 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8225 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8226 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8227 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8228 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8229 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8230 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8231 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8232 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8233 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8234 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8235 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8236 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8237 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8238 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8239 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8240 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8241 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8242 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8243 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8244 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8245 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8246 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8247 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8248 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8249 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8250 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8251 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8252 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8253 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8254 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8255 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8256 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8257 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8258 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8259 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8260 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8261 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8262 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8263 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8264 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8265 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8266 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8267 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8268 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8269 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8270 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8271 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8272 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8273 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8274 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8275 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8276 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8277 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8278 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8279 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8280 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8281 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8282 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8283 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8284 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8285 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8286 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8287 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8288 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8289 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8290 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8291 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8292 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8293 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8294 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8295 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8296 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8297 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8298 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8299 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8300 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8301 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8302 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8303 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8304 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8305 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8306 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8307 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8308 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8309 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8310 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8311 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8312 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8313 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8314 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8315 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8316 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8317 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8318 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8319 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8320 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8321 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8322 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8323 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8324 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8325 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8326 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8327 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8328 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8329 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8330 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8331 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8332 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8333 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8334 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8335 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8336 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8337 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8338 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8339 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8340 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8341 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8342 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8343 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8344 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8345 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8346 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8347 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8348 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8349 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8350 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8351 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8352 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8353 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8354 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8355 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8356 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8357 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8358 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8359 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8360 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8361 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8362 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8363 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8364 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8365 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8366 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8367 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8368 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8369 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8370 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8371 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8372 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8373 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8374 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8375 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8376 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8377 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8378 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8379 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8380 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8381 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8382 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8383 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8384 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8385 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8386 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8387 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8388 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8389 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8390 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8391 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8392 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8393 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8394 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8395 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8396 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8397 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8398 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8399 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8400 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8401 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8402 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8403 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8404 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8405 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8406 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8407 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8408 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8409 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8410 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8411 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8412 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8413 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8414 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8415 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8416 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8417 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8418 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8419 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8420 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8421 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8422 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8423 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8424 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8425 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8426 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8427 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8428 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8429 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8430 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8431 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8432 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8433 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8434 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8435 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8436 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8437 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8438 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8439 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8440 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8441 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8442 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8443 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8444 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8445 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8446 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8447 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8448 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8449 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8450 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8451 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8452 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8453 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8454 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8455 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8456 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8457 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8458 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8459 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8460 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8461 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8462 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8463 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8464 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8465 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8466 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8467 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8468 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8469 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8470 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8471 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8472 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8473 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8474 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8475 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8476 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8477 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8478 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8479 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8480 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8481 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8482 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8483 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8484 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8485 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8486 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8487 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8488 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8489 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8490 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8491 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8492 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8493 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8494 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8495 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8496 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8497 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8498 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8499 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8500 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8501 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8502 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8503 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8504 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8505 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8506 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8507 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8508 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8509 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8510 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8511 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8512 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8513 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8514 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8515 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8516 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8517 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8518 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8519 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8520 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8521 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8522 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8523 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8524 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8525 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8526 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8527 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8528 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8529 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8530 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8531 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8532 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8533 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8534 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8535 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8536 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8537 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8538 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8539 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8540 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8541 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8542 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8543 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8544 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8545 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8546 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8547 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8548 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8549 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8550 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8551 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8552 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8553 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8554 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8555 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8556 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8557 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8558 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8559 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8560 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8561 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8562 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8563 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8564 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8565 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8566 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8567 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8568 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8569 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8570 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8571 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8572 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8573 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8574 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8575 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8576 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8577 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8578 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8579 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8580 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8581 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8582 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8583 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8584 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8585 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8586 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8587 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8588 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8589 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8590 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8591 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8592 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8593 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8594 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8595 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8596 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8597 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8598 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8599 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8600 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8601 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8602 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8603 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8604 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8605 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8606 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8607 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8608 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8609 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8610 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8611 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8612 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8613 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8614 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8615 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8616 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8617 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8618 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8619 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8620 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8621 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8622 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8623 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8624 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8625 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8626 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8627 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8628 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8629 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8630 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8631 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8632 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8633 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8634 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8635 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8636 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8637 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8638 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8639 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8640 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8641 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8642 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8643 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8644 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8645 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8646 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8647 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8648 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8649 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8650 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8651 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8652 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8653 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8654 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8655 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8656 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8657 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8658 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8659 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8660 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8661 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8662 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8663 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8664 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8665 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8666 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8667 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8668 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8669 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8670 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8671 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8672 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8673 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8674 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8675 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8676 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8677 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8678 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8679 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8680 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8681 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8682 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8683 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8684 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8685 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8686 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8687 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8688 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8689 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8690 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8691 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8692 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8693 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8694 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8695 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8696 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8697 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8698 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8699 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8700 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8701 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8702 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8703 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8704 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8705 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8706 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8707 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8708 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8709 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8710 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8711 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8712 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8713 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8714 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8715 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8716 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8717 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8718 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8719 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8720 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8721 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8722 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8723 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8724 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8725 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8726 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8727 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8728 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8729 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8730 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8731 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8732 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8733 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8734 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8735 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8736 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8737 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8738 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8739 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8740 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8741 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8742 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8743 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8744 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8745 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8746 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8747 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8748 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8749 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8750 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8751 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8752 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8753 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8754 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8755 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8756 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8757 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8758 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8759 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8760 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8761 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8762 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8763 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8764 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8765 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8766 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8767 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8768 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8769 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8770 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8771 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8772 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8773 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8774 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8775 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8776 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8777 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8778 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8779 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8780 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8781 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8782 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8783 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8784 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8785 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8786 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8787 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8788 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8789 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8790 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8791 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8792 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8793 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8794 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8795 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8796 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8797 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8798 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8799 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8800 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8801 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8802 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8803 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8804 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8805 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8806 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8807 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8808 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8809 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8810 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8811 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8812 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8813 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8814 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8815 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8816 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8817 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8818 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8819 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8820 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8821 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8822 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8823 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8824 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8825 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8826 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8827 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8828 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8829 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8830 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8831 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8832 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8833 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8834 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8835 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8836 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8837 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8838 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8839 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8840 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8841 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8842 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8843 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8844 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8845 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8846 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8847 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8848 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8849 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8850 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8851 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8852 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8853 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8854 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8855 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8856 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8857 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8858 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8859 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8860 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8861 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8862 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8863 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8864 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8865 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8866 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8867 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8868 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8869 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8870 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8871 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8872 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8873 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8874 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8875 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8876 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8877 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8878 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8879 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8880 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8881 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8882 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8883 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8884 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8885 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8886 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8887 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8888 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8889 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8890 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8891 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8892 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8893 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8894 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8895 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8896 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8897 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8898 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8899 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8900 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8901 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8902 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8903 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8904 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8905 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8906 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8907 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8908 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8909 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8910 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8911 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8912 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8913 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8914 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8915 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8916 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8917 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8918 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8919 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8920 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8921 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8922 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8923 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8924 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8925 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8926 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8927 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8928 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8929 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8930 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8931 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8932 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8933 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8934 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8935 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8936 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8937 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8938 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8939 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8940 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8941 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8942 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8943 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8944 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8945 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8946 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8947 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8948 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8949 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8950 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8951 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8952 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8953 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8954 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8955 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8956 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8957 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8958 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8959 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8960 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8961 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8962 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8963 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8964 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8965 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8966 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8967 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8968 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8969 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8970 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8971 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8972 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8973 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8974 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8975 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8976 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8977 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8978 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8979 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8980 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8981 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8982 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8983 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8984 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8985 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8986 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8987 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8988 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8989 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8990 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8991 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8992 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8993 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8994 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8995 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8996 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8997 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8998 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		8999 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9000 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9001 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9002 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9003 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9004 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9005 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9006 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9007 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9008 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9009 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9010 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9011 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9012 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9013 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9014 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9015 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9016 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9017 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9018 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9019 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9020 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9021 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9022 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9023 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9024 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9025 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9026 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9027 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9028 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9029 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9030 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9031 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9032 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9033 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9034 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9035 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9036 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9037 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9038 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9039 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9040 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9041 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9042 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9043 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9044 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9045 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9046 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9047 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9048 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9049 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9050 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9051 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9052 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9053 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9054 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9055 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9056 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9057 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9058 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9059 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9060 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9061 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9062 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9063 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9064 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9065 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9066 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9067 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9068 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9069 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9070 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9071 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9072 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9073 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9074 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9075 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9076 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9077 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9078 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9079 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9080 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9081 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9082 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9083 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9084 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9085 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9086 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		9087 =>	x"000063FF", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"
	);


--			***** COLOR PALLETE *****




begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;